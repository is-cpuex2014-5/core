library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

library UNISIM;
use UNISIM.VComponents.all;

-- CPUEV2(HW09) より
entity top is
  Port (MCLK1   : in    STD_LOGIC;
         RS_TX  : out   STD_LOGIC;
         XGA    : out   STD_LOGIC;
         XE1    : out   STD_LOGIC;
         E2A    : out   STD_LOGIC;
         XE3    : out   STD_LOGIC;
         XZCKE  : out   STD_LOGIC;
         ADVA   : out   STD_LOGIC;
         XLBO   : out   STD_LOGIC;
         ZZA    : out   STD_LOGIC;
         XFT    : out   STD_LOGIC;
         ZCLKMA : out   STD_LOGIC_VECTOR (1 downto 0);
         ZD     : inout STD_LOGIC_VECTOR (31 downto 0);
         ZDP    : inout STD_LOGIC_VECTOR (3 downto 0);
         ZA     : inout STD_LOGIC_VECTOR (19 downto 0);
         IOA    :       STD_LOGIC_VECTOR (126 downto 0);
         XZBE   : inout STD_LOGIC_VECTOR (3 downto 0);
         XWA    : out   STD_LOGIC;
         XRST   : in    STD_LOGIC;
         RS_RX  : in    STD_LOGIC);
end top;

architecture cpu_top of top is
  signal clk,iclk : std_logic;
  --testbench signal
  component core Port (
    clk                   : in  std_logic;
    execute_ok            : in  std_logic;
    ostate                : out std_logic_vector(7 downto 0);
    sram_go               : out std_logic;
    sram_inst_type        : out std_logic;
    sram_addr             : out std_logic_vector(19 downto 0);
    sram_read             : in  std_logic_vector(31 downto 0);
    sram_write            : out std_logic_vector(31 downto 0);
    debug_otpt            : out std_logic_vector(7 downto 0);
    debug_otpt_signal     : out std_logic;
    waitwrite_from_parent : in  std_logic_vector(19 downto 0);
    read_signal           : out std_logic
  );
  end component;
  component sram Port (
    clk            : in    std_logic;
    SRXGA          : out   STD_LOGIC;
    SRXE1          : out   STD_LOGIC;
    SRE2A          : out   STD_LOGIC;
    SRXE3          : out   STD_LOGIC;
    SRXZCKE        : out   STD_LOGIC;
    SRADVA         : out   STD_LOGIC;
    SRXLBO         : out   STD_LOGIC;
    SRZZA          : out   STD_LOGIC;
    SRXFT          : out   STD_LOGIC;
    SRZCLKMA       : out   STD_LOGIC_VECTOR (1 downto 0);
    SRZD           : inout STD_LOGIC_VECTOR (31 downto 0);
    SRZDP          : inout STD_LOGIC_VECTOR (3 downto 0);
    SRZA           : inout STD_LOGIC_VECTOR (19 downto 0);
    SRIOA          :       STD_LOGIC_VECTOR (126 downto 0);
    SRXZBE         : inout STD_LOGIC_VECTOR (3 downto 0);
    SRXWA          : out   STD_LOGIC;
    SRXRST         : in    STD_LOGIC;
    sram_go        : in    std_logic;
    sram_busy      : out   std_logic;
    sram_inst_type : in    std_logic;
    sram_read      : out   std_logic_vector(31 downto 0);
    sram_write     : in    std_logic_vector(31 downto 0);
    sram_addr      : in    std_logic_vector(19 downto 0)
  );
  end component;
  component u232c
    generic (wtime: std_logic_vector(15 downto 0) := x"1ADB");
    Port (
      clk      : in  std_logic;
      data_reg : in  std_logic_vector(7 downto 0);
      go       : in  std_logic;
      busy     : out std_logic;
      tx       : out std_logic
    );
  end component;
  component inputc
    Port (
      clk         : in  std_logic;
      execute_ok  : out std_logic;
      debug_read  : out std_logic_vector(7 downto 0);
      write_value : out std_logic_vector(31 downto 0);
      write_addr  : out std_logic_vector(19 downto 0);
      write_ok    : out std_logic;
      rx          : in  std_logic
    );
  end component;
  component write_buff is
    generic (
      buff_size : integer range 0 to 65535);
    port (
      clk      : in  std_logic;
      data_in  : in  std_logic_vector (7 downto 0);
      go_in    : in  std_logic;
      busy_in  : in  std_logic;
      data_out : out std_logic_vector (7 downto 0);
      go_out   : out std_logic;
      busy_out : out std_logic);
  end component write_buff;

  signal exok : std_logic := '0';
  signal exok_from_read : std_logic := '0';
  signal top_state : std_logic := '0';
  signal hogge : std_logic_vector(7 downto 0);
  signal debug_otpt : std_logic_vector(7 downto 0);
  signal debug_otpt_signal : std_logic;
  signal debug_otpt_inputc : std_logic_vector(7 downto 0);
  signal u232c_data_reg : std_logic_vector(7 downto 0);
  signal u232c_go : std_logic := '0';
  signal u232c_busy : std_logic;
  signal inputc_write_value : std_logic_vector(31 downto 0);
  signal inputc_write_addr : std_logic_vector(19 downto 0);
  signal inputc_write_ok : std_logic;
  signal core_sram_go : std_logic;
  signal core_sram_inst_type : std_logic; --0: read 1: write
  signal core_sram_read : std_logic_vector(31 downto 0);
  signal core_sram_write : std_logic_vector(31 downto 0);
  signal core_sram_addr : std_logic_vector(19 downto 0);
  signal sram_go : std_logic;
  signal sram_busy : std_logic;
  signal sram_inst_type : std_logic; --0: read 1: write
  signal sram_read : std_logic_vector(31 downto 0);
  signal sram_write : std_logic_vector(31 downto 0);
  signal sram_addr : std_logic_vector(19 downto 0);
  signal sigcount : std_logic_vector(3 downto 0) := x"0";
  signal debug_saved_value : std_logic_vector(31 downto 0);
  signal first_state_sram_input_id : std_logic_vector(19 downto 0) := x"00000";
  signal first_state_write_wait : std_logic_vector(7 downto 0) := x"00";
  signal waitwrite_to_core : std_logic_vector(19 downto 0) := x"00000";
  -- wait one clock to wait u232c's busy
  signal debug_waitoneclock : std_logic := '0';
  signal read_signal : std_logic;
  signal read_inst_addr : std_logic_vector(19 downto 0) := x"55554";
  signal sram_read_transfer_mode : std_logic := '0'; -- 0: normal  1: read_signal_ver
  signal read_counter : std_logic_vector(1 downto 0) := "00";
  signal read_counter_old : std_logic_vector(1 downto 0) := "00";
  signal write_buff_busy : std_logic := '0';
begin
  -- HW 実験当時の top より
  ib: IBUFG port map (
    i => MCLK1,
    o => iclk
    );
  bg: BUFG port map (
    i => iclk,
    o => clk
    );
  rs232c : u232c generic map (wtime => x"1ADB")
  Port map (
    clk      => clk,
    data_reg => u232c_data_reg,
    go       => u232c_go,
    busy     => u232c_busy,
    tx       => rs_tx
    );
  with_inputc : inputc Port map (
    clk         => clk,
    execute_ok  => exok_from_read,
    debug_read  => debug_otpt_inputc,
    write_value => inputc_write_value,
    write_addr  => inputc_write_addr,
    write_ok    => inputc_write_ok,
    rx          => rs_rx
    );
  core_send: core Port map (
    clk                   => clk,
    execute_ok            => exok,
    ostate                => hogge,
    sram_go               => core_sram_go,
    sram_inst_type        => core_sram_inst_type,
    sram_read             => core_sram_read,
    sram_write            => core_sram_write,
    sram_addr             => core_sram_addr,
    debug_otpt            => debug_otpt,
    debug_otpt_signal     => debug_otpt_signal,
    waitwrite_from_parent => waitwrite_to_core,
    read_signal           => read_signal
    );
  withsram: sram Port map (
    clk            => clk,
    SRXGA          => XGA,
    SRXE1          => XE1,
    SRE2A          => E2A,
    SRXE3          => XE3,
    SRXZCKE        => XZCKE,
    SRADVA         => ADVA,
    SRXLBO         => XLBO,
    SRZZA          => ZZA,
    SRXFT          => XFT,
    SRZCLKMA       => ZCLKMA,
    SRZD           => ZD,
    SRZDP          => ZDP,
    SRZA           => ZA,
    SRIOA          => IOA,
    SRXZBE         => XZBE,
    SRXWA          => XWA,
    SRXRST         => XRST,
    sram_go        => sram_go,
    sram_busy      => sram_busy,
    sram_inst_type => sram_inst_type,
    sram_read      => sram_read,
    sram_write     => sram_write,
    sram_addr      => sram_addr
    );
  with_write_buff: write_buff
    generic map (
      buff_size => 256)
    port map (
      clk      => clk,
      data_in  => debug_otpt,
      go_in    => debug_otpt_signal,
      busy_in  => u232c_busy,
      data_out => u232c_data_reg,
      go_out   => u232c_go,
      busy_out => write_buff_busy);

  cpu_top_main : process
  begin
    if rising_edge(clk) then
      if write_buff_busy = '0' then
        waitwrite_to_core <= x"00000";
      else
        waitwrite_to_core <= x"C0C0A";
      end if;
      if top_state = '0' then
        --Input Wait
        if exok_from_read = '1' then
          exok      <= '1';
          top_state <= '1';
        end if;
        if sram_busy = '0' then
          if inputc_write_ok = '1' then
            sram_go           <= '1';
            --write
            sram_inst_type    <= '1';
            sram_addr         <= inputc_write_addr;
            sram_write        <= inputc_write_value;
            debug_saved_value <= inputc_write_value;
            sigcount          <= x"8";
          else
            sram_go <= '0';
          end if;
        else
          sram_go <= '0';
        end if;
      end if;
      if top_state = '1' then
        if sram_read_transfer_mode = '1' then
          -- read 命令
          if read_counter_old = 0 then
            core_sram_read <= x"000000" & sram_read(7 downto 0);
          end if;
          if read_counter_old = 1 then
            core_sram_read <= x"000000" & sram_read(15 downto 8);
          end if;
          if read_counter_old = 2 then
            core_sram_read <= x"000000" & sram_read(23 downto 16);
          end if;
          if read_counter_old = 3 then
            core_sram_read <= x"000000" & sram_read(31 downto 24);
          end if;
        else
          -- 垂れ流し
          core_sram_read <= sram_read;
        end if;
        if read_signal = '1' then
          if sram_busy = '0' then
            sram_go        <= '1';
            sram_inst_type <= '0';
            sram_addr      <= read_inst_addr;
            if read_counter = 3 then
              read_inst_addr <= read_inst_addr - 1;
            end if;
            read_counter_old        <= read_counter;
            read_counter            <= read_counter + 1;
            sram_read_transfer_mode <= '1';
          end if;
        else
          if sram_busy = '0' then
            if core_sram_go = '1' then
              sram_go <= '1';
              if core_sram_inst_type = '0' then
                --read
                sram_inst_type          <= '0';
                sram_addr               <= core_sram_addr;
                sram_read_transfer_mode <= '0';
              else
                --write
                sram_inst_type <= '1';
                sram_addr      <= core_sram_addr;
                sram_write     <= core_sram_write;
              end if;
            else
              sram_go <= '0';
            end if;
          else
            sram_go <= '0';
          end if;
        end if;
      end if;
    end if;
  end process;
end cpu_top;

