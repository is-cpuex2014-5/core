library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

library UNISIM;
use UNISIM.VComponents.all;

-- CPUEV2(HW09) より
entity top is
  Port ( MCLK1 : in  STD_LOGIC;
         RS_TX : out  STD_LOGIC;
         XGA : out STD_LOGIC;
         XE1 : out STD_LOGIC;
         E2A : out STD_LOGIC;
         XE3 : out STD_LOGIC;
         XZCKE : out STD_LOGIC;
         ADVA : out STD_LOGIC;
         XLBO : out STD_LOGIC;
         ZZA : out STD_LOGIC;
         XFT : out STD_LOGIC;
         ZCLKMA : out STD_LOGIC_VECTOR (1 downto 0);
         ZD : inout STD_LOGIC_VECTOR (31 downto 0);
         ZDP : inout STD_LOGIC_VECTOR (3 downto 0);
         ZA : inout STD_LOGIC_VECTOR (19 downto 0);
         IOA : STD_LOGIC_VECTOR (126 downto 0);
         XZBE : inout STD_LOGIC_VECTOR (3 downto 0);
         XWA : out STD_LOGIC;
         XRST : in STD_LOGIC;
         RS_RX : in STD_LOGIC
        );
end top;

architecture cpu_top of top is
  signal clk,iclk : std_logic;
  --testbench signal
  component core Port (
    clk: in std_logic;
    execute_ok: in std_logic;
    ostate: out std_logic_vector(7 downto 0);
    sram_go : out std_logic;
    sram_inst_type : out std_logic;
    sram_addr : out std_logic_vector(19 downto 0);
    sram_read : in std_logic_vector(31 downto 0);
    sram_write : out std_logic_vector(31 downto 0);
    debug_otpt: out std_logic_vector(31 downto 0);
    debug_otpt_code: out std_logic_vector(2 downto 0);
    debug_otpt_signal: out std_logic;
    waitwrite_from_parent : in std_logic_vector(19 downto 0)
  );
  end component;
  component sram Port (
    clk: in std_logic;
    SRXGA : out STD_LOGIC;
    SRXE1 : out STD_LOGIC;
    SRE2A : out STD_LOGIC;
    SRXE3 : out STD_LOGIC;
    SRXZCKE : out STD_LOGIC;
    SRADVA : out STD_LOGIC;
    SRXLBO : out STD_LOGIC;
    SRZZA : out STD_LOGIC;
    SRXFT : out STD_LOGIC;
    SRZCLKMA : out STD_LOGIC_VECTOR (1 downto 0);
    SRZD : inout STD_LOGIC_VECTOR (31 downto 0);
    SRZDP : inout STD_LOGIC_VECTOR (3 downto 0);
    SRZA : inout STD_LOGIC_VECTOR (19 downto 0);
    SRIOA : STD_LOGIC_VECTOR (126 downto 0);
    SRXZBE : inout STD_LOGIC_VECTOR (3 downto 0);
    SRXWA : out STD_LOGIC;
    SRXRST : in STD_LOGIC;
    sram_go : in std_logic;
    sram_busy : out std_logic;
    sram_inst_type : in std_logic;
    sram_read : out std_logic_vector(31 downto 0);
    sram_write : in std_logic_vector(31 downto 0);
    sram_addr : in std_logic_vector(19 downto 0)
  );
  end component;
  component u232c
    generic (wtime: std_logic_vector(15 downto 0) := x"1ADB");
    Port (
      clk : in std_logic;
      data_reg : in std_logic_vector(31 downto 0);
      showtype : in std_logic_vector(2 downto 0);
      go : in std_logic;
      busy : out std_logic;
      tx : out std_logic
    );
  end component;
  component inputc
    Port (
      clk : in std_logic;
      execute_ok : out std_logic;
      debug_read : out std_logic_vector(7 downto 0);
      write_value : out std_logic_vector(31 downto 0);
      write_addr : out std_logic_vector(19 downto 0);
      write_ok : out std_logic;
      rx : in std_logic
    );
  end component;
  signal exok : std_logic := '0';
  signal exok_from_read : std_logic;
  signal top_state : std_logic_vector(2 downto 0) := "000";
  signal hogge : std_logic_vector(7 downto 0);
  signal debug_otpt : std_logic_vector(31 downto 0);
  signal debug_otpt_code : std_logic_vector(2 downto 0);
  signal debug_otpt_signal : std_logic;
  signal debug_otpt_inputc : std_logic_vector(7 downto 0);
  signal u232c_data_reg : std_logic_vector(31 downto 0);
  signal u232c_showtype : std_logic_vector(2 downto 0);
  signal u232c_go : std_logic;
  signal u232c_busy : std_logic;
  signal inputc_write_value : std_logic_vector(31 downto 0);
  signal inputc_write_addr : std_logic_vector(19 downto 0);
  signal inputc_write_ok : std_logic;
  signal core_sram_go : std_logic;
  signal core_sram_inst_type : std_logic; --0: read 1: write
  signal core_sram_read : std_logic_vector(31 downto 0);
  signal core_sram_write : std_logic_vector(31 downto 0);
  signal core_sram_addr : std_logic_vector(19 downto 0);
  signal sram_go : std_logic;
  signal sram_busy : std_logic;
  signal sram_inst_type : std_logic; --0: read 1: write
  signal sram_read : std_logic_vector(31 downto 0);
  signal sram_write : std_logic_vector(31 downto 0);
  signal sram_addr : std_logic_vector(19 downto 0);
  signal sigcount : std_logic_vector(3 downto 0) := x"0";
  signal debug_saved_value : std_logic_vector(31 downto 0);
  signal first_state_sram_input_id : std_logic_vector(19 downto 0) := x"00000";
  signal first_state_write_wait : std_logic_vector(7 downto 0) := x"00";
  signal waitwrite_to_core : std_logic_vector(19 downto 0) := x"00000";
  -- wait one clock to wait u232c's busy
  signal debug_waitoneclock : std_logic := '0';
begin
  -- HW 実験当時の top より
  ib: IBUFG port map (
    i => MCLK1,
    o => iclk
    );
  bg: BUFG port map (
    i => iclk,
    o => clk
    );
  rs232c : u232c generic map (wtime => x"1ADB")
  Port map (
    clk => clk,
    data_reg => u232c_data_reg,
    showtype => u232c_showtype,
    go => u232c_go,
    busy => u232c_busy,
    tx => rs_tx
    );
  with_inputc : inputc Port map (
    clk => clk,
    execute_ok => exok_from_read,
    debug_read => debug_otpt_inputc,
    write_value => inputc_write_value,
    write_addr => inputc_write_addr,
    write_ok => inputc_write_ok,
    rx => rs_rx
    );
  core_send: core Port map (
    clk => clk,
    execute_ok => exok,
    ostate => hogge,
    sram_go => core_sram_go,
    sram_inst_type => core_sram_inst_type,
    sram_read => core_sram_read,
    sram_write => core_sram_write,
    sram_addr => core_sram_addr,
    debug_otpt => debug_otpt,
    debug_otpt_code => debug_otpt_code,
    debug_otpt_signal => debug_otpt_signal,
    waitwrite_from_parent => waitwrite_to_core
    );
  withsram: sram Port map (
    clk => clk,
    SRXGA => XGA,
    SRXE1 => XE1,
    SRE2A => E2A,
    SRXE3 => XE3,
    SRXZCKE => XZCKE,
    SRADVA => ADVA,
    SRXLBO => XLBO,
    SRZZA => ZZA,
    SRXFT => XFT,
    SRZCLKMA => ZCLKMA,
    SRZD => ZD,
    SRZDP => ZDP,
    SRZA => ZA,
    SRIOA => IOA,
    SRXZBE => XZBE,
    SRXWA => XWA,
    SRXRST => XRST,
    sram_go => sram_go,
    sram_busy => sram_busy,
    sram_inst_type => sram_inst_type,
    sram_read => sram_read,
    sram_write => sram_write,
    sram_addr => sram_addr
    );
  cpu_top_main : process
  begin
    if rising_edge(clk) then
      if u232c_busy = '0' then
        waitwrite_to_core <= x"00000";
      else
        waitwrite_to_core <= x"C0C0A";
      end if;
      if top_state = "000" then
        -- write inst phase
        if (first_state_write_wait = 0) then
        -- write in addr
          if (first_state_sram_input_id<15522) then
            if sram_busy = '0' then
              sram_go <= '1';
              sram_inst_type <= '1';
              first_state_write_wait <= x"FF";
              sram_addr <= first_state_sram_input_id;
if first_state_sram_input_id = 0 then
	sram_write <= x"8200F250";
end if;
if first_state_sram_input_id = 1 then
	sram_write <= x"43000000";
end if;
if first_state_sram_input_id = 2 then
	sram_write <= x"BDCCCCCD";
end if;
if first_state_sram_input_id = 3 then
	sram_write <= x"3F666666";
end if;
if first_state_sram_input_id = 4 then
	sram_write <= x"3E4CCCCD";
end if;
if first_state_sram_input_id = 5 then
	sram_write <= x"C3160000";
end if;
if first_state_sram_input_id = 6 then
	sram_write <= x"43160000";
end if;
if first_state_sram_input_id = 7 then
	sram_write <= x"3DCCCCCD";
end if;
if first_state_sram_input_id = 8 then
	sram_write <= x"C0000000";
end if;
if first_state_sram_input_id = 9 then
	sram_write <= x"43800000";
end if;
if first_state_sram_input_id = 10 then
	sram_write <= x"4CBEBC20";
end if;
if first_state_sram_input_id = 11 then
	sram_write <= x"4E6E6B28";
end if;
if first_state_sram_input_id = 12 then
	sram_write <= x"41A00000";
end if;
if first_state_sram_input_id = 13 then
	sram_write <= x"3D4CCCCD";
end if;
if first_state_sram_input_id = 14 then
	sram_write <= x"3E800000";
end if;
if first_state_sram_input_id = 15 then
	sram_write <= x"41200000";
end if;
if first_state_sram_input_id = 16 then
	sram_write <= x"3E99999A";
end if;
if first_state_sram_input_id = 17 then
	sram_write <= x"437F0000";
end if;
if first_state_sram_input_id = 18 then
	sram_write <= x"3E19999A";
end if;
if first_state_sram_input_id = 19 then
	sram_write <= x"41700000";
end if;
if first_state_sram_input_id = 20 then
	sram_write <= x"40490FDC";
end if;
if first_state_sram_input_id = 21 then
	sram_write <= x"41F00000";
end if;
if first_state_sram_input_id = 22 then
	sram_write <= x"3C75989E";
end if;
if first_state_sram_input_id = 23 then
	sram_write <= x"3F6DA101";
end if;
if first_state_sram_input_id = 24 then
	sram_write <= x"3C8F53C5";
end if;
if first_state_sram_input_id = 25 then
	sram_write <= x"3E0E9468";
end if;
if first_state_sram_input_id = 26 then
	sram_write <= x"3CF30835";
end if;
if first_state_sram_input_id = 27 then
	sram_write <= x"38D1B717";
end if;
if first_state_sram_input_id = 28 then
	sram_write <= x"BDCCCCCD";
end if;
if first_state_sram_input_id = 29 then
	sram_write <= x"3C23D70A";
end if;
if first_state_sram_input_id = 30 then
	sram_write <= x"BE4CCCCD";
end if;
if first_state_sram_input_id = 31 then
	sram_write <= x"BF800000";
end if;
if first_state_sram_input_id = 32 then
	sram_write <= x"40000000";
end if;
if first_state_sram_input_id = 33 then
	sram_write <= x"C3480000";
end if;
if first_state_sram_input_id = 34 then
	sram_write <= x"43480000";
end if;
if first_state_sram_input_id = 35 then
	sram_write <= x"3C8EF998";
end if;
if first_state_sram_input_id = 36 then
	sram_write <= x"C0C90FDA";
end if;
if first_state_sram_input_id = 37 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 38 then
	sram_write <= x"40C90FDA";
end if;
if first_state_sram_input_id = 39 then
	sram_write <= x"3AB39192";
end if;
if first_state_sram_input_id = 40 then
	sram_write <= x"3D2AA7DF";
end if;
if first_state_sram_input_id = 41 then
	sram_write <= x"3F000000";
end if;
if first_state_sram_input_id = 42 then
	sram_write <= x"3F800000";
end if;
if first_state_sram_input_id = 43 then
	sram_write <= x"394D8559";
end if;
if first_state_sram_input_id = 44 then
	sram_write <= x"3C088723";
end if;
if first_state_sram_input_id = 45 then
	sram_write <= x"3E2AAAC1";
end if;
if first_state_sram_input_id = 46 then
	sram_write <= x"3F490FD8";
end if;
if first_state_sram_input_id = 47 then
	sram_write <= x"3FC90FD8";
end if;
if first_state_sram_input_id = 48 then
	sram_write <= x"40490FDC";
end if;
if first_state_sram_input_id = 49 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 50 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 51 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 52 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 53 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 54 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 55 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 56 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 57 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 58 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 59 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 60 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 61 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 62 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 63 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 64 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 65 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 66 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 67 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 68 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 69 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 70 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 71 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 72 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 73 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 74 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 75 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 76 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 77 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 78 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 79 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 80 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 81 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 82 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 83 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 84 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 85 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 86 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 87 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 88 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 89 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 90 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 91 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 92 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 93 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 94 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 95 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 96 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 97 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 98 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 99 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 100 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 101 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 102 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 103 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 104 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 105 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 106 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 107 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 108 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 109 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 110 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 111 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 112 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 113 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 114 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 115 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 116 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 117 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 118 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 119 then
	sram_write <= x"437F0000";
end if;
if first_state_sram_input_id = 120 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 121 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 122 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 123 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 124 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 125 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 126 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 127 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 128 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 129 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 130 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 131 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 132 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 133 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 134 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 135 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 136 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 137 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 138 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 139 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 140 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 141 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 142 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 143 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 144 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 145 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 146 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 147 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 148 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 149 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 150 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 151 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 152 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 153 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 154 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 155 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 156 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 157 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 158 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 159 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 160 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 161 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 162 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 163 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 164 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 165 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 166 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 167 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 168 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 169 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 170 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 171 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 172 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 173 then
	sram_write <= x"4E6E6B28";
end if;
if first_state_sram_input_id = 174 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 175 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 176 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 177 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 178 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 179 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 180 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 181 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 182 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 183 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 184 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 185 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 186 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 187 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 188 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 189 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 190 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 191 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 192 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 193 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 194 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 195 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 196 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 197 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 198 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 199 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 200 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 201 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 202 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 203 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 204 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 205 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 206 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 207 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 208 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 209 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 210 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 211 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 212 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 213 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 214 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 215 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 216 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 217 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 218 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 219 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 220 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 221 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 222 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 223 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 224 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 225 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 226 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 227 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 228 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 229 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 230 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 231 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 232 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 233 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 234 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 235 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 236 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 237 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 238 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 239 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 240 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 241 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 242 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 243 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 244 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 245 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 246 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 247 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 248 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 249 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 250 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 251 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 252 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 253 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 254 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 255 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 256 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 257 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 258 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 259 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 260 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 261 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 262 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 263 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 264 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 265 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 266 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 267 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 268 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 269 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 270 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 271 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 272 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 273 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 274 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 275 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 276 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 277 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 278 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 279 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 280 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 281 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 282 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 283 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 284 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 285 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 286 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 287 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 288 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 289 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 290 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 291 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 292 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 293 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 294 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 295 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 296 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 297 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 298 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 299 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 300 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 301 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 302 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 303 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 304 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 305 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 306 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 307 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 308 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 309 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 310 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 311 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 312 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 313 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 314 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 315 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 316 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 317 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 318 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 319 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 320 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 321 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 322 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 323 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 324 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 325 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 326 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 327 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 328 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 329 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 330 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 331 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 332 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 333 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 334 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 335 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 336 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 337 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 338 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 339 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 340 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 341 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 342 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 343 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 344 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 345 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 346 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 347 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 348 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 349 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 350 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 351 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 352 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 353 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 354 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 355 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 356 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 357 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 358 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 359 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 360 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 361 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 362 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 363 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 364 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 365 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 366 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 367 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 368 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 369 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 370 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 371 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 372 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 373 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 374 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 375 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 376 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 377 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 378 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 379 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 380 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 381 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 382 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 383 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 384 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 385 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 386 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 387 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 388 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 389 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 390 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 391 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 392 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 393 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 394 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 395 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 396 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 397 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 398 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 399 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 400 then
	sram_write <= x"00000000";
end if;
if first_state_sram_input_id = 401 then
	sram_write <= x"028000EC";
end if;
if first_state_sram_input_id = 402 then
	sram_write <= x"02A000C8";
end if;
if first_state_sram_input_id = 403 then
	sram_write <= x"06C00001";
end if;
if first_state_sram_input_id = 404 then
	sram_write <= x"0220000B";
end if;
if first_state_sram_input_id = 405 then
	sram_write <= x"02400000";
end if;
if first_state_sram_input_id = 406 then
	sram_write <= x"03DC0004";
end if;
if first_state_sram_input_id = 407 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 408 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 409 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 410 then
	sram_write <= x"07DC0004";
end if;
if first_state_sram_input_id = 411 then
	sram_write <= x"0048A000";
end if;
if first_state_sram_input_id = 412 then
	sram_write <= x"C4240000";
end if;
if first_state_sram_input_id = 413 then
	sram_write <= x"06880004";
end if;
if first_state_sram_input_id = 414 then
	sram_write <= x"86C80650";
end if;
if first_state_sram_input_id = 415 then
	sram_write <= x"028000C4";
end if;
if first_state_sram_input_id = 416 then
	sram_write <= x"02A001E0";
end if;
if first_state_sram_input_id = 417 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 418 then
	sram_write <= x"0240FFFF";
end if;
if first_state_sram_input_id = 419 then
	sram_write <= x"03DC0004";
end if;
if first_state_sram_input_id = 420 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 421 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 422 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 423 then
	sram_write <= x"07DC0004";
end if;
if first_state_sram_input_id = 424 then
	sram_write <= x"0048A000";
end if;
if first_state_sram_input_id = 425 then
	sram_write <= x"C4240000";
end if;
if first_state_sram_input_id = 426 then
	sram_write <= x"06880004";
end if;
if first_state_sram_input_id = 427 then
	sram_write <= x"86C80684";
end if;
if first_state_sram_input_id = 428 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 429 then
	sram_write <= x"0240FFFF";
end if;
if first_state_sram_input_id = 430 then
	sram_write <= x"03DC0004";
end if;
if first_state_sram_input_id = 431 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 432 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 433 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 434 then
	sram_write <= x"07DC0004";
end if;
if first_state_sram_input_id = 435 then
	sram_write <= x"00420000";
end if;
if first_state_sram_input_id = 436 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 437 then
	sram_write <= x"03DC0004";
end if;
if first_state_sram_input_id = 438 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 439 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 440 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 441 then
	sram_write <= x"07DC0004";
end if;
if first_state_sram_input_id = 442 then
	sram_write <= x"C42002A8";
end if;
if first_state_sram_input_id = 443 then
	sram_write <= x"02A00368";
end if;
if first_state_sram_input_id = 444 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 445 then
	sram_write <= x"02400000";
end if;
if first_state_sram_input_id = 446 then
	sram_write <= x"03DC0004";
end if;
if first_state_sram_input_id = 447 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 448 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 449 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 450 then
	sram_write <= x"07DC0004";
end if;
if first_state_sram_input_id = 451 then
	sram_write <= x"C42A0000";
end if;
if first_state_sram_input_id = 452 then
	sram_write <= x"0220003C";
end if;
if first_state_sram_input_id = 453 then
	sram_write <= x"03DC0004";
end if;
if first_state_sram_input_id = 454 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 455 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 456 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 457 then
	sram_write <= x"07DC0004";
end if;
if first_state_sram_input_id = 458 then
	sram_write <= x"C42A0004";
end if;
if first_state_sram_input_id = 459 then
	sram_write <= x"028002CC";
end if;
if first_state_sram_input_id = 460 then
	sram_write <= x"02A00370";
end if;
if first_state_sram_input_id = 461 then
	sram_write <= x"02200002";
end if;
if first_state_sram_input_id = 462 then
	sram_write <= x"03DC0004";
end if;
if first_state_sram_input_id = 463 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 464 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 465 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 466 then
	sram_write <= x"07DC0004";
end if;
if first_state_sram_input_id = 467 then
	sram_write <= x"00E20000";
end if;
if first_state_sram_input_id = 468 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 469 then
	sram_write <= x"02400000";
end if;
if first_state_sram_input_id = 470 then
	sram_write <= x"03DC0004";
end if;
if first_state_sram_input_id = 471 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 472 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 473 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 474 then
	sram_write <= x"07DC0004";
end if;
if first_state_sram_input_id = 475 then
	sram_write <= x"C4E20004";
end if;
if first_state_sram_input_id = 476 then
	sram_write <= x"0048A000";
end if;
if first_state_sram_input_id = 477 then
	sram_write <= x"C4240000";
end if;
if first_state_sram_input_id = 478 then
	sram_write <= x"06880004";
end if;
if first_state_sram_input_id = 479 then
	sram_write <= x"86C80734";
end if;
if first_state_sram_input_id = 480 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 481 then
	sram_write <= x"E0200000";
end if;
if first_state_sram_input_id = 482 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 483 then
	sram_write <= x"E2200000";
end if;
if first_state_sram_input_id = 484 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 485 then
	sram_write <= x"E0200000";
end if;
if first_state_sram_input_id = 486 then
	sram_write <= x"E0400000";
end if;
if first_state_sram_input_id = 487 then
	sram_write <= x"E0600000";
end if;
if first_state_sram_input_id = 488 then
	sram_write <= x"E0800000";
end if;
if first_state_sram_input_id = 489 then
	sram_write <= x"22221820";
end if;
if first_state_sram_input_id = 490 then
	sram_write <= x"22441020";
end if;
if first_state_sram_input_id = 491 then
	sram_write <= x"22660820";
end if;
if first_state_sram_input_id = 492 then
	sram_write <= x"00224000";
end if;
if first_state_sram_input_id = 493 then
	sram_write <= x"00226000";
end if;
if first_state_sram_input_id = 494 then
	sram_write <= x"00228000";
end if;
if first_state_sram_input_id = 495 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 496 then
	sram_write <= x"E0200000";
end if;
if first_state_sram_input_id = 497 then
	sram_write <= x"E0400000";
end if;
if first_state_sram_input_id = 498 then
	sram_write <= x"E0600000";
end if;
if first_state_sram_input_id = 499 then
	sram_write <= x"E0800000";
end if;
if first_state_sram_input_id = 500 then
	sram_write <= x"22221820";
end if;
if first_state_sram_input_id = 501 then
	sram_write <= x"22441020";
end if;
if first_state_sram_input_id = 502 then
	sram_write <= x"22660820";
end if;
if first_state_sram_input_id = 503 then
	sram_write <= x"00224000";
end if;
if first_state_sram_input_id = 504 then
	sram_write <= x"00226000";
end if;
if first_state_sram_input_id = 505 then
	sram_write <= x"00228000";
end if;
if first_state_sram_input_id = 506 then
	sram_write <= x"C43C0004";
end if;
if first_state_sram_input_id = 507 then
	sram_write <= x"C83C0004";
end if;
if first_state_sram_input_id = 508 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 509 then
	sram_write <= x"CC3C0004";
end if;
if first_state_sram_input_id = 510 then
	sram_write <= x"C03C0004";
end if;
if first_state_sram_input_id = 511 then
	sram_write <= x"228218A0";
end if;
if first_state_sram_input_id = 512 then
	sram_write <= x"226210A0";
end if;
if first_state_sram_input_id = 513 then
	sram_write <= x"224208A0";
end if;
if first_state_sram_input_id = 514 then
	sram_write <= x"E2800000";
end if;
if first_state_sram_input_id = 515 then
	sram_write <= x"E2600000";
end if;
if first_state_sram_input_id = 516 then
	sram_write <= x"E2400000";
end if;
if first_state_sram_input_id = 517 then
	sram_write <= x"E2200000";
end if;
if first_state_sram_input_id = 518 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 519 then
	sram_write <= x"007A0000";
end if;
if first_state_sram_input_id = 520 then
	sram_write <= x"82200834";
end if;
if first_state_sram_input_id = 521 then
	sram_write <= x"C45A0000";
end if;
if first_state_sram_input_id = 522 then
	sram_write <= x"06220001";
end if;
if first_state_sram_input_id = 523 then
	sram_write <= x"03BA0004";
end if;
if first_state_sram_input_id = 524 then
	sram_write <= x"82000820";
end if;
if first_state_sram_input_id = 525 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 526 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 527 then
	sram_write <= x"50220000";
end if;
if first_state_sram_input_id = 528 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 529 then
	sram_write <= x"60220000";
end if;
if first_state_sram_input_id = 530 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 531 then
	sram_write <= x"C84000C0";
end if;
if first_state_sram_input_id = 532 then
	sram_write <= x"C86000BC";
end if;
if first_state_sram_input_id = 533 then
	sram_write <= x"C88000B8";
end if;
if first_state_sram_input_id = 534 then
	sram_write <= x"C43C0000";
end if;
if first_state_sram_input_id = 535 then
	sram_write <= x"8E240A10";
end if;
if first_state_sram_input_id = 536 then
	sram_write <= x"44224000";
end if;
if first_state_sram_input_id = 537 then
	sram_write <= x"04402000";
end if;
if first_state_sram_input_id = 538 then
	sram_write <= x"C45C0004";
end if;
if first_state_sram_input_id = 539 then
	sram_write <= x"8E240898";
end if;
if first_state_sram_input_id = 540 then
	sram_write <= x"44224000";
end if;
if first_state_sram_input_id = 541 then
	sram_write <= x"04604000";
end if;
if first_state_sram_input_id = 542 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 543 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 544 then
	sram_write <= x"03DC0010";
end if;
if first_state_sram_input_id = 545 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 546 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 547 then
	sram_write <= x"8200084C";
end if;
if first_state_sram_input_id = 548 then
	sram_write <= x"07DC0010";
end if;
if first_state_sram_input_id = 549 then
	sram_write <= x"820009F8";
end if;
if first_state_sram_input_id = 550 then
	sram_write <= x"8E26094C";
end if;
if first_state_sram_input_id = 551 then
	sram_write <= x"8E8208F8";
end if;
if first_state_sram_input_id = 552 then
	sram_write <= x"C84000B4";
end if;
if first_state_sram_input_id = 553 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 554 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 555 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 556 then
	sram_write <= x"44424000";
end if;
if first_state_sram_input_id = 557 then
	sram_write <= x"C86000B0";
end if;
if first_state_sram_input_id = 558 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 559 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 560 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 561 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 562 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 563 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 564 then
	sram_write <= x"C86000AC";
end if;
if first_state_sram_input_id = 565 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 566 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 567 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 568 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 569 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 570 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 571 then
	sram_write <= x"48262000";
end if;
if first_state_sram_input_id = 572 then
	sram_write <= x"44242000";
end if;
if first_state_sram_input_id = 573 then
	sram_write <= x"82000948";
end if;
if first_state_sram_input_id = 574 then
	sram_write <= x"44262000";
end if;
if first_state_sram_input_id = 575 then
	sram_write <= x"C84000A8";
end if;
if first_state_sram_input_id = 576 then
	sram_write <= x"C86000A4";
end if;
if first_state_sram_input_id = 577 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 578 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 579 then
	sram_write <= x"44446000";
end if;
if first_state_sram_input_id = 580 then
	sram_write <= x"C86000A0";
end if;
if first_state_sram_input_id = 581 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 582 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 583 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 584 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 585 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 586 then
	sram_write <= x"C860009C";
end if;
if first_state_sram_input_id = 587 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 588 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 589 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 590 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 591 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 592 then
	sram_write <= x"48262000";
end if;
if first_state_sram_input_id = 593 then
	sram_write <= x"44242000";
end if;
if first_state_sram_input_id = 594 then
	sram_write <= x"820009F8";
end if;
if first_state_sram_input_id = 595 then
	sram_write <= x"8E8209A8";
end if;
if first_state_sram_input_id = 596 then
	sram_write <= x"C84000B4";
end if;
if first_state_sram_input_id = 597 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 598 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 599 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 600 then
	sram_write <= x"44424000";
end if;
if first_state_sram_input_id = 601 then
	sram_write <= x"C86000B0";
end if;
if first_state_sram_input_id = 602 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 603 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 604 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 605 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 606 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 607 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 608 then
	sram_write <= x"C86000AC";
end if;
if first_state_sram_input_id = 609 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 610 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 611 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 612 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 613 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 614 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 615 then
	sram_write <= x"48262000";
end if;
if first_state_sram_input_id = 616 then
	sram_write <= x"44242000";
end if;
if first_state_sram_input_id = 617 then
	sram_write <= x"820009F8";
end if;
if first_state_sram_input_id = 618 then
	sram_write <= x"44262000";
end if;
if first_state_sram_input_id = 619 then
	sram_write <= x"C84000A8";
end if;
if first_state_sram_input_id = 620 then
	sram_write <= x"C86000A4";
end if;
if first_state_sram_input_id = 621 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 622 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 623 then
	sram_write <= x"44446000";
end if;
if first_state_sram_input_id = 624 then
	sram_write <= x"C86000A0";
end if;
if first_state_sram_input_id = 625 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 626 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 627 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 628 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 629 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 630 then
	sram_write <= x"C860009C";
end if;
if first_state_sram_input_id = 631 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 632 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 633 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 634 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 635 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 636 then
	sram_write <= x"48262000";
end if;
if first_state_sram_input_id = 637 then
	sram_write <= x"44242000";
end if;
if first_state_sram_input_id = 638 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 639 then
	sram_write <= x"C05C0004";
end if;
if first_state_sram_input_id = 640 then
	sram_write <= x"82420A08";
end if;
if first_state_sram_input_id = 641 then
	sram_write <= x"82000A0C";
end if;
if first_state_sram_input_id = 642 then
	sram_write <= x"44202000";
end if;
if first_state_sram_input_id = 643 then
	sram_write <= x"82000B70";
end if;
if first_state_sram_input_id = 644 then
	sram_write <= x"8E260AC4";
end if;
if first_state_sram_input_id = 645 then
	sram_write <= x"8E820A70";
end if;
if first_state_sram_input_id = 646 then
	sram_write <= x"C84000B4";
end if;
if first_state_sram_input_id = 647 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 648 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 649 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 650 then
	sram_write <= x"44424000";
end if;
if first_state_sram_input_id = 651 then
	sram_write <= x"C86000B0";
end if;
if first_state_sram_input_id = 652 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 653 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 654 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 655 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 656 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 657 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 658 then
	sram_write <= x"C86000AC";
end if;
if first_state_sram_input_id = 659 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 660 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 661 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 662 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 663 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 664 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 665 then
	sram_write <= x"48262000";
end if;
if first_state_sram_input_id = 666 then
	sram_write <= x"44242000";
end if;
if first_state_sram_input_id = 667 then
	sram_write <= x"82000AC0";
end if;
if first_state_sram_input_id = 668 then
	sram_write <= x"44262000";
end if;
if first_state_sram_input_id = 669 then
	sram_write <= x"C84000A8";
end if;
if first_state_sram_input_id = 670 then
	sram_write <= x"C86000A4";
end if;
if first_state_sram_input_id = 671 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 672 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 673 then
	sram_write <= x"44446000";
end if;
if first_state_sram_input_id = 674 then
	sram_write <= x"C86000A0";
end if;
if first_state_sram_input_id = 675 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 676 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 677 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 678 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 679 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 680 then
	sram_write <= x"C860009C";
end if;
if first_state_sram_input_id = 681 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 682 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 683 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 684 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 685 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 686 then
	sram_write <= x"48262000";
end if;
if first_state_sram_input_id = 687 then
	sram_write <= x"44242000";
end if;
if first_state_sram_input_id = 688 then
	sram_write <= x"82000B70";
end if;
if first_state_sram_input_id = 689 then
	sram_write <= x"8E820B20";
end if;
if first_state_sram_input_id = 690 then
	sram_write <= x"C84000B4";
end if;
if first_state_sram_input_id = 691 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 692 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 693 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 694 then
	sram_write <= x"44424000";
end if;
if first_state_sram_input_id = 695 then
	sram_write <= x"C86000B0";
end if;
if first_state_sram_input_id = 696 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 697 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 698 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 699 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 700 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 701 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 702 then
	sram_write <= x"C86000AC";
end if;
if first_state_sram_input_id = 703 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 704 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 705 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 706 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 707 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 708 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 709 then
	sram_write <= x"48262000";
end if;
if first_state_sram_input_id = 710 then
	sram_write <= x"44242000";
end if;
if first_state_sram_input_id = 711 then
	sram_write <= x"82000B70";
end if;
if first_state_sram_input_id = 712 then
	sram_write <= x"44262000";
end if;
if first_state_sram_input_id = 713 then
	sram_write <= x"C84000A8";
end if;
if first_state_sram_input_id = 714 then
	sram_write <= x"C86000A4";
end if;
if first_state_sram_input_id = 715 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 716 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 717 then
	sram_write <= x"44446000";
end if;
if first_state_sram_input_id = 718 then
	sram_write <= x"C86000A0";
end if;
if first_state_sram_input_id = 719 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 720 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 721 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 722 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 723 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 724 then
	sram_write <= x"C860009C";
end if;
if first_state_sram_input_id = 725 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 726 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 727 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 728 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 729 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 730 then
	sram_write <= x"48262000";
end if;
if first_state_sram_input_id = 731 then
	sram_write <= x"44242000";
end if;
if first_state_sram_input_id = 732 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 733 then
	sram_write <= x"C05C0000";
end if;
if first_state_sram_input_id = 734 then
	sram_write <= x"82420B80";
end if;
if first_state_sram_input_id = 735 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 736 then
	sram_write <= x"44202000";
end if;
if first_state_sram_input_id = 737 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 738 then
	sram_write <= x"C84000C0";
end if;
if first_state_sram_input_id = 739 then
	sram_write <= x"C86000BC";
end if;
if first_state_sram_input_id = 740 then
	sram_write <= x"C88000B8";
end if;
if first_state_sram_input_id = 741 then
	sram_write <= x"C43C0000";
end if;
if first_state_sram_input_id = 742 then
	sram_write <= x"8E240D4C";
end if;
if first_state_sram_input_id = 743 then
	sram_write <= x"44224000";
end if;
if first_state_sram_input_id = 744 then
	sram_write <= x"04402000";
end if;
if first_state_sram_input_id = 745 then
	sram_write <= x"C45C0004";
end if;
if first_state_sram_input_id = 746 then
	sram_write <= x"8E240BD4";
end if;
if first_state_sram_input_id = 747 then
	sram_write <= x"44224000";
end if;
if first_state_sram_input_id = 748 then
	sram_write <= x"04604000";
end if;
if first_state_sram_input_id = 749 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 750 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 751 then
	sram_write <= x"03DC0010";
end if;
if first_state_sram_input_id = 752 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 753 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 754 then
	sram_write <= x"8200084C";
end if;
if first_state_sram_input_id = 755 then
	sram_write <= x"07DC0010";
end if;
if first_state_sram_input_id = 756 then
	sram_write <= x"82000D34";
end if;
if first_state_sram_input_id = 757 then
	sram_write <= x"8E260C88";
end if;
if first_state_sram_input_id = 758 then
	sram_write <= x"8E820C34";
end if;
if first_state_sram_input_id = 759 then
	sram_write <= x"C84000B4";
end if;
if first_state_sram_input_id = 760 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 761 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 762 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 763 then
	sram_write <= x"44424000";
end if;
if first_state_sram_input_id = 764 then
	sram_write <= x"C86000B0";
end if;
if first_state_sram_input_id = 765 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 766 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 767 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 768 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 769 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 770 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 771 then
	sram_write <= x"C86000AC";
end if;
if first_state_sram_input_id = 772 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 773 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 774 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 775 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 776 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 777 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 778 then
	sram_write <= x"48262000";
end if;
if first_state_sram_input_id = 779 then
	sram_write <= x"44242000";
end if;
if first_state_sram_input_id = 780 then
	sram_write <= x"82000C84";
end if;
if first_state_sram_input_id = 781 then
	sram_write <= x"44262000";
end if;
if first_state_sram_input_id = 782 then
	sram_write <= x"C84000A8";
end if;
if first_state_sram_input_id = 783 then
	sram_write <= x"C86000A4";
end if;
if first_state_sram_input_id = 784 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 785 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 786 then
	sram_write <= x"44446000";
end if;
if first_state_sram_input_id = 787 then
	sram_write <= x"C86000A0";
end if;
if first_state_sram_input_id = 788 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 789 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 790 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 791 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 792 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 793 then
	sram_write <= x"C860009C";
end if;
if first_state_sram_input_id = 794 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 795 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 796 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 797 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 798 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 799 then
	sram_write <= x"48262000";
end if;
if first_state_sram_input_id = 800 then
	sram_write <= x"44242000";
end if;
if first_state_sram_input_id = 801 then
	sram_write <= x"82000D34";
end if;
if first_state_sram_input_id = 802 then
	sram_write <= x"8E820CE4";
end if;
if first_state_sram_input_id = 803 then
	sram_write <= x"C84000B4";
end if;
if first_state_sram_input_id = 804 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 805 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 806 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 807 then
	sram_write <= x"44424000";
end if;
if first_state_sram_input_id = 808 then
	sram_write <= x"C86000B0";
end if;
if first_state_sram_input_id = 809 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 810 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 811 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 812 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 813 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 814 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 815 then
	sram_write <= x"C86000AC";
end if;
if first_state_sram_input_id = 816 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 817 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 818 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 819 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 820 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 821 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 822 then
	sram_write <= x"48262000";
end if;
if first_state_sram_input_id = 823 then
	sram_write <= x"44242000";
end if;
if first_state_sram_input_id = 824 then
	sram_write <= x"82000D34";
end if;
if first_state_sram_input_id = 825 then
	sram_write <= x"44262000";
end if;
if first_state_sram_input_id = 826 then
	sram_write <= x"C84000A8";
end if;
if first_state_sram_input_id = 827 then
	sram_write <= x"C86000A4";
end if;
if first_state_sram_input_id = 828 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 829 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 830 then
	sram_write <= x"44446000";
end if;
if first_state_sram_input_id = 831 then
	sram_write <= x"C86000A0";
end if;
if first_state_sram_input_id = 832 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 833 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 834 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 835 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 836 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 837 then
	sram_write <= x"C860009C";
end if;
if first_state_sram_input_id = 838 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 839 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 840 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 841 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 842 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 843 then
	sram_write <= x"48262000";
end if;
if first_state_sram_input_id = 844 then
	sram_write <= x"44242000";
end if;
if first_state_sram_input_id = 845 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 846 then
	sram_write <= x"C05C0004";
end if;
if first_state_sram_input_id = 847 then
	sram_write <= x"82420D44";
end if;
if first_state_sram_input_id = 848 then
	sram_write <= x"82000D48";
end if;
if first_state_sram_input_id = 849 then
	sram_write <= x"44202000";
end if;
if first_state_sram_input_id = 850 then
	sram_write <= x"82000EAC";
end if;
if first_state_sram_input_id = 851 then
	sram_write <= x"8E260E00";
end if;
if first_state_sram_input_id = 852 then
	sram_write <= x"8E820DA4";
end if;
if first_state_sram_input_id = 853 then
	sram_write <= x"C84000A8";
end if;
if first_state_sram_input_id = 854 then
	sram_write <= x"C86000A4";
end if;
if first_state_sram_input_id = 855 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 856 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 857 then
	sram_write <= x"44446000";
end if;
if first_state_sram_input_id = 858 then
	sram_write <= x"C86000A0";
end if;
if first_state_sram_input_id = 859 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 860 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 861 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 862 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 863 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 864 then
	sram_write <= x"C860009C";
end if;
if first_state_sram_input_id = 865 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 866 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 867 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 868 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 869 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 870 then
	sram_write <= x"48262000";
end if;
if first_state_sram_input_id = 871 then
	sram_write <= x"44242000";
end if;
if first_state_sram_input_id = 872 then
	sram_write <= x"82000DFC";
end if;
if first_state_sram_input_id = 873 then
	sram_write <= x"44262000";
end if;
if first_state_sram_input_id = 874 then
	sram_write <= x"C84000B4";
end if;
if first_state_sram_input_id = 875 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 876 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 877 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 878 then
	sram_write <= x"44424000";
end if;
if first_state_sram_input_id = 879 then
	sram_write <= x"C86000B0";
end if;
if first_state_sram_input_id = 880 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 881 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 882 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 883 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 884 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 885 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 886 then
	sram_write <= x"C86000AC";
end if;
if first_state_sram_input_id = 887 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 888 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 889 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 890 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 891 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 892 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 893 then
	sram_write <= x"48262000";
end if;
if first_state_sram_input_id = 894 then
	sram_write <= x"44242000";
end if;
if first_state_sram_input_id = 895 then
	sram_write <= x"82000EAC";
end if;
if first_state_sram_input_id = 896 then
	sram_write <= x"8E820E54";
end if;
if first_state_sram_input_id = 897 then
	sram_write <= x"C84000A8";
end if;
if first_state_sram_input_id = 898 then
	sram_write <= x"C86000A4";
end if;
if first_state_sram_input_id = 899 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 900 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 901 then
	sram_write <= x"44446000";
end if;
if first_state_sram_input_id = 902 then
	sram_write <= x"C86000A0";
end if;
if first_state_sram_input_id = 903 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 904 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 905 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 906 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 907 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 908 then
	sram_write <= x"C860009C";
end if;
if first_state_sram_input_id = 909 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 910 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 911 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 912 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 913 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 914 then
	sram_write <= x"48262000";
end if;
if first_state_sram_input_id = 915 then
	sram_write <= x"44242000";
end if;
if first_state_sram_input_id = 916 then
	sram_write <= x"82000EAC";
end if;
if first_state_sram_input_id = 917 then
	sram_write <= x"44262000";
end if;
if first_state_sram_input_id = 918 then
	sram_write <= x"C84000B4";
end if;
if first_state_sram_input_id = 919 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 920 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 921 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 922 then
	sram_write <= x"44424000";
end if;
if first_state_sram_input_id = 923 then
	sram_write <= x"C86000B0";
end if;
if first_state_sram_input_id = 924 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 925 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 926 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 927 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 928 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 929 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 930 then
	sram_write <= x"C86000AC";
end if;
if first_state_sram_input_id = 931 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 932 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 933 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 934 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 935 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 936 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 937 then
	sram_write <= x"48262000";
end if;
if first_state_sram_input_id = 938 then
	sram_write <= x"44242000";
end if;
if first_state_sram_input_id = 939 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 940 then
	sram_write <= x"C05C0000";
end if;
if first_state_sram_input_id = 941 then
	sram_write <= x"82420EBC";
end if;
if first_state_sram_input_id = 942 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 943 then
	sram_write <= x"44202000";
end if;
if first_state_sram_input_id = 944 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 945 then
	sram_write <= x"C8400098";
end if;
if first_state_sram_input_id = 946 then
	sram_write <= x"8E240F00";
end if;
if first_state_sram_input_id = 947 then
	sram_write <= x"44224000";
end if;
if first_state_sram_input_id = 948 then
	sram_write <= x"8E240EDC";
end if;
if first_state_sram_input_id = 949 then
	sram_write <= x"44224000";
end if;
if first_state_sram_input_id = 950 then
	sram_write <= x"82000EC4";
end if;
if first_state_sram_input_id = 951 then
	sram_write <= x"8E020EF8";
end if;
if first_state_sram_input_id = 952 then
	sram_write <= x"C8600090";
end if;
if first_state_sram_input_id = 953 then
	sram_write <= x"8E620EF0";
end if;
if first_state_sram_input_id = 954 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 955 then
	sram_write <= x"82000EC4";
end if;
if first_state_sram_input_id = 956 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 957 then
	sram_write <= x"8200084C";
end if;
if first_state_sram_input_id = 958 then
	sram_write <= x"0220FFFF";
end if;
if first_state_sram_input_id = 959 then
	sram_write <= x"8200084C";
end if;
if first_state_sram_input_id = 960 then
	sram_write <= x"8E0210D8";
end if;
if first_state_sram_input_id = 961 then
	sram_write <= x"C8600090";
end if;
if first_state_sram_input_id = 962 then
	sram_write <= x"8E620F3C";
end if;
if first_state_sram_input_id = 963 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 964 then
	sram_write <= x"8E240F1C";
end if;
if first_state_sram_input_id = 965 then
	sram_write <= x"44224000";
end if;
if first_state_sram_input_id = 966 then
	sram_write <= x"82000EC4";
end if;
if first_state_sram_input_id = 967 then
	sram_write <= x"8E020F34";
end if;
if first_state_sram_input_id = 968 then
	sram_write <= x"8E620F2C";
end if;
if first_state_sram_input_id = 969 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 970 then
	sram_write <= x"82000EC4";
end if;
if first_state_sram_input_id = 971 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 972 then
	sram_write <= x"8200084C";
end if;
if first_state_sram_input_id = 973 then
	sram_write <= x"0220FFFF";
end if;
if first_state_sram_input_id = 974 then
	sram_write <= x"8200084C";
end if;
if first_state_sram_input_id = 975 then
	sram_write <= x"C84000C0";
end if;
if first_state_sram_input_id = 976 then
	sram_write <= x"C86000BC";
end if;
if first_state_sram_input_id = 977 then
	sram_write <= x"C88000B8";
end if;
if first_state_sram_input_id = 978 then
	sram_write <= x"8E240F70";
end if;
if first_state_sram_input_id = 979 then
	sram_write <= x"44224000";
end if;
if first_state_sram_input_id = 980 then
	sram_write <= x"0220FFFF";
end if;
if first_state_sram_input_id = 981 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 982 then
	sram_write <= x"03DC0008";
end if;
if first_state_sram_input_id = 983 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 984 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 985 then
	sram_write <= x"8200084C";
end if;
if first_state_sram_input_id = 986 then
	sram_write <= x"07DC0008";
end if;
if first_state_sram_input_id = 987 then
	sram_write <= x"820010D0";
end if;
if first_state_sram_input_id = 988 then
	sram_write <= x"8E261024";
end if;
if first_state_sram_input_id = 989 then
	sram_write <= x"8E820FD0";
end if;
if first_state_sram_input_id = 990 then
	sram_write <= x"C84000B4";
end if;
if first_state_sram_input_id = 991 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 992 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 993 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 994 then
	sram_write <= x"44424000";
end if;
if first_state_sram_input_id = 995 then
	sram_write <= x"C86000B0";
end if;
if first_state_sram_input_id = 996 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 997 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 998 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 999 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1000 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1001 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 1002 then
	sram_write <= x"C86000AC";
end if;
if first_state_sram_input_id = 1003 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1004 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1005 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1006 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1007 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1008 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1009 then
	sram_write <= x"48262000";
end if;
if first_state_sram_input_id = 1010 then
	sram_write <= x"44242000";
end if;
if first_state_sram_input_id = 1011 then
	sram_write <= x"82001020";
end if;
if first_state_sram_input_id = 1012 then
	sram_write <= x"44262000";
end if;
if first_state_sram_input_id = 1013 then
	sram_write <= x"C84000A8";
end if;
if first_state_sram_input_id = 1014 then
	sram_write <= x"C86000A4";
end if;
if first_state_sram_input_id = 1015 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1016 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1017 then
	sram_write <= x"44446000";
end if;
if first_state_sram_input_id = 1018 then
	sram_write <= x"C86000A0";
end if;
if first_state_sram_input_id = 1019 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1020 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1021 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1022 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1023 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 1024 then
	sram_write <= x"C860009C";
end if;
if first_state_sram_input_id = 1025 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1026 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1027 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1028 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1029 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1030 then
	sram_write <= x"48262000";
end if;
if first_state_sram_input_id = 1031 then
	sram_write <= x"44242000";
end if;
if first_state_sram_input_id = 1032 then
	sram_write <= x"820010D0";
end if;
if first_state_sram_input_id = 1033 then
	sram_write <= x"8E821080";
end if;
if first_state_sram_input_id = 1034 then
	sram_write <= x"C84000B4";
end if;
if first_state_sram_input_id = 1035 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 1036 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 1037 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 1038 then
	sram_write <= x"44424000";
end if;
if first_state_sram_input_id = 1039 then
	sram_write <= x"C86000B0";
end if;
if first_state_sram_input_id = 1040 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1041 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1042 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1043 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1044 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1045 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 1046 then
	sram_write <= x"C86000AC";
end if;
if first_state_sram_input_id = 1047 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1048 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1049 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1050 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1051 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1052 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1053 then
	sram_write <= x"48262000";
end if;
if first_state_sram_input_id = 1054 then
	sram_write <= x"44242000";
end if;
if first_state_sram_input_id = 1055 then
	sram_write <= x"820010D0";
end if;
if first_state_sram_input_id = 1056 then
	sram_write <= x"44262000";
end if;
if first_state_sram_input_id = 1057 then
	sram_write <= x"C84000A8";
end if;
if first_state_sram_input_id = 1058 then
	sram_write <= x"C86000A4";
end if;
if first_state_sram_input_id = 1059 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1060 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1061 then
	sram_write <= x"44446000";
end if;
if first_state_sram_input_id = 1062 then
	sram_write <= x"C86000A0";
end if;
if first_state_sram_input_id = 1063 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1064 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1065 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1066 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1067 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 1068 then
	sram_write <= x"C860009C";
end if;
if first_state_sram_input_id = 1069 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1070 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1071 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1072 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1073 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1074 then
	sram_write <= x"48262000";
end if;
if first_state_sram_input_id = 1075 then
	sram_write <= x"44242000";
end if;
if first_state_sram_input_id = 1076 then
	sram_write <= x"44202000";
end if;
if first_state_sram_input_id = 1077 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 1078 then
	sram_write <= x"C84000C0";
end if;
if first_state_sram_input_id = 1079 then
	sram_write <= x"C86000BC";
end if;
if first_state_sram_input_id = 1080 then
	sram_write <= x"C88000B8";
end if;
if first_state_sram_input_id = 1081 then
	sram_write <= x"8E24110C";
end if;
if first_state_sram_input_id = 1082 then
	sram_write <= x"44224000";
end if;
if first_state_sram_input_id = 1083 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 1084 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1085 then
	sram_write <= x"03DC0008";
end if;
if first_state_sram_input_id = 1086 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1087 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1088 then
	sram_write <= x"8200084C";
end if;
if first_state_sram_input_id = 1089 then
	sram_write <= x"07DC0008";
end if;
if first_state_sram_input_id = 1090 then
	sram_write <= x"8200126C";
end if;
if first_state_sram_input_id = 1091 then
	sram_write <= x"8E2611C0";
end if;
if first_state_sram_input_id = 1092 then
	sram_write <= x"8E82116C";
end if;
if first_state_sram_input_id = 1093 then
	sram_write <= x"C84000B4";
end if;
if first_state_sram_input_id = 1094 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 1095 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 1096 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 1097 then
	sram_write <= x"44424000";
end if;
if first_state_sram_input_id = 1098 then
	sram_write <= x"C86000B0";
end if;
if first_state_sram_input_id = 1099 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1100 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1101 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1102 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1103 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1104 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 1105 then
	sram_write <= x"C86000AC";
end if;
if first_state_sram_input_id = 1106 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1107 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1108 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1109 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1110 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1111 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1112 then
	sram_write <= x"48262000";
end if;
if first_state_sram_input_id = 1113 then
	sram_write <= x"44242000";
end if;
if first_state_sram_input_id = 1114 then
	sram_write <= x"820011BC";
end if;
if first_state_sram_input_id = 1115 then
	sram_write <= x"44262000";
end if;
if first_state_sram_input_id = 1116 then
	sram_write <= x"C84000A8";
end if;
if first_state_sram_input_id = 1117 then
	sram_write <= x"C86000A4";
end if;
if first_state_sram_input_id = 1118 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1119 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1120 then
	sram_write <= x"44446000";
end if;
if first_state_sram_input_id = 1121 then
	sram_write <= x"C86000A0";
end if;
if first_state_sram_input_id = 1122 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1123 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1124 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1125 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1126 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 1127 then
	sram_write <= x"C860009C";
end if;
if first_state_sram_input_id = 1128 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1129 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1130 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1131 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1132 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1133 then
	sram_write <= x"48262000";
end if;
if first_state_sram_input_id = 1134 then
	sram_write <= x"44242000";
end if;
if first_state_sram_input_id = 1135 then
	sram_write <= x"8200126C";
end if;
if first_state_sram_input_id = 1136 then
	sram_write <= x"8E82121C";
end if;
if first_state_sram_input_id = 1137 then
	sram_write <= x"C84000B4";
end if;
if first_state_sram_input_id = 1138 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 1139 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 1140 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 1141 then
	sram_write <= x"44424000";
end if;
if first_state_sram_input_id = 1142 then
	sram_write <= x"C86000B0";
end if;
if first_state_sram_input_id = 1143 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1144 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1145 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1146 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1147 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1148 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 1149 then
	sram_write <= x"C86000AC";
end if;
if first_state_sram_input_id = 1150 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1151 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1152 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1153 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1154 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1155 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1156 then
	sram_write <= x"48262000";
end if;
if first_state_sram_input_id = 1157 then
	sram_write <= x"44242000";
end if;
if first_state_sram_input_id = 1158 then
	sram_write <= x"8200126C";
end if;
if first_state_sram_input_id = 1159 then
	sram_write <= x"44262000";
end if;
if first_state_sram_input_id = 1160 then
	sram_write <= x"C84000A8";
end if;
if first_state_sram_input_id = 1161 then
	sram_write <= x"C86000A4";
end if;
if first_state_sram_input_id = 1162 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1163 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1164 then
	sram_write <= x"44446000";
end if;
if first_state_sram_input_id = 1165 then
	sram_write <= x"C86000A0";
end if;
if first_state_sram_input_id = 1166 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1167 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1168 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1169 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1170 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 1171 then
	sram_write <= x"C860009C";
end if;
if first_state_sram_input_id = 1172 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1173 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1174 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1175 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1176 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1177 then
	sram_write <= x"48262000";
end if;
if first_state_sram_input_id = 1178 then
	sram_write <= x"44242000";
end if;
if first_state_sram_input_id = 1179 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 1180 then
	sram_write <= x"C8400098";
end if;
if first_state_sram_input_id = 1181 then
	sram_write <= x"8E2412AC";
end if;
if first_state_sram_input_id = 1182 then
	sram_write <= x"44224000";
end if;
if first_state_sram_input_id = 1183 then
	sram_write <= x"8E241288";
end if;
if first_state_sram_input_id = 1184 then
	sram_write <= x"44224000";
end if;
if first_state_sram_input_id = 1185 then
	sram_write <= x"82001270";
end if;
if first_state_sram_input_id = 1186 then
	sram_write <= x"8E0212A4";
end if;
if first_state_sram_input_id = 1187 then
	sram_write <= x"C8600090";
end if;
if first_state_sram_input_id = 1188 then
	sram_write <= x"8E62129C";
end if;
if first_state_sram_input_id = 1189 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 1190 then
	sram_write <= x"82001270";
end if;
if first_state_sram_input_id = 1191 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 1192 then
	sram_write <= x"82000B88";
end if;
if first_state_sram_input_id = 1193 then
	sram_write <= x"0220FFFF";
end if;
if first_state_sram_input_id = 1194 then
	sram_write <= x"82000B88";
end if;
if first_state_sram_input_id = 1195 then
	sram_write <= x"8E021484";
end if;
if first_state_sram_input_id = 1196 then
	sram_write <= x"C8600090";
end if;
if first_state_sram_input_id = 1197 then
	sram_write <= x"8E6212E8";
end if;
if first_state_sram_input_id = 1198 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 1199 then
	sram_write <= x"8E2412C8";
end if;
if first_state_sram_input_id = 1200 then
	sram_write <= x"44224000";
end if;
if first_state_sram_input_id = 1201 then
	sram_write <= x"82001270";
end if;
if first_state_sram_input_id = 1202 then
	sram_write <= x"8E0212E0";
end if;
if first_state_sram_input_id = 1203 then
	sram_write <= x"8E6212D8";
end if;
if first_state_sram_input_id = 1204 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 1205 then
	sram_write <= x"82001270";
end if;
if first_state_sram_input_id = 1206 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 1207 then
	sram_write <= x"82000B88";
end if;
if first_state_sram_input_id = 1208 then
	sram_write <= x"0220FFFF";
end if;
if first_state_sram_input_id = 1209 then
	sram_write <= x"82000B88";
end if;
if first_state_sram_input_id = 1210 then
	sram_write <= x"C84000C0";
end if;
if first_state_sram_input_id = 1211 then
	sram_write <= x"C86000BC";
end if;
if first_state_sram_input_id = 1212 then
	sram_write <= x"C88000B8";
end if;
if first_state_sram_input_id = 1213 then
	sram_write <= x"8E24131C";
end if;
if first_state_sram_input_id = 1214 then
	sram_write <= x"44224000";
end if;
if first_state_sram_input_id = 1215 then
	sram_write <= x"0220FFFF";
end if;
if first_state_sram_input_id = 1216 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1217 then
	sram_write <= x"03DC0008";
end if;
if first_state_sram_input_id = 1218 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1219 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1220 then
	sram_write <= x"8200084C";
end if;
if first_state_sram_input_id = 1221 then
	sram_write <= x"07DC0008";
end if;
if first_state_sram_input_id = 1222 then
	sram_write <= x"8200147C";
end if;
if first_state_sram_input_id = 1223 then
	sram_write <= x"8E2613D0";
end if;
if first_state_sram_input_id = 1224 then
	sram_write <= x"8E821374";
end if;
if first_state_sram_input_id = 1225 then
	sram_write <= x"C84000A8";
end if;
if first_state_sram_input_id = 1226 then
	sram_write <= x"C86000A4";
end if;
if first_state_sram_input_id = 1227 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1228 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1229 then
	sram_write <= x"44446000";
end if;
if first_state_sram_input_id = 1230 then
	sram_write <= x"C86000A0";
end if;
if first_state_sram_input_id = 1231 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1232 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1233 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1234 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1235 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 1236 then
	sram_write <= x"C860009C";
end if;
if first_state_sram_input_id = 1237 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1238 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1239 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1240 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1241 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1242 then
	sram_write <= x"48262000";
end if;
if first_state_sram_input_id = 1243 then
	sram_write <= x"44242000";
end if;
if first_state_sram_input_id = 1244 then
	sram_write <= x"820013CC";
end if;
if first_state_sram_input_id = 1245 then
	sram_write <= x"44262000";
end if;
if first_state_sram_input_id = 1246 then
	sram_write <= x"C84000B4";
end if;
if first_state_sram_input_id = 1247 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 1248 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 1249 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 1250 then
	sram_write <= x"44424000";
end if;
if first_state_sram_input_id = 1251 then
	sram_write <= x"C86000B0";
end if;
if first_state_sram_input_id = 1252 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1253 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1254 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1255 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1256 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1257 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 1258 then
	sram_write <= x"C86000AC";
end if;
if first_state_sram_input_id = 1259 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1260 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1261 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1262 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1263 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1264 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1265 then
	sram_write <= x"48262000";
end if;
if first_state_sram_input_id = 1266 then
	sram_write <= x"44242000";
end if;
if first_state_sram_input_id = 1267 then
	sram_write <= x"8200147C";
end if;
if first_state_sram_input_id = 1268 then
	sram_write <= x"8E821424";
end if;
if first_state_sram_input_id = 1269 then
	sram_write <= x"C84000A8";
end if;
if first_state_sram_input_id = 1270 then
	sram_write <= x"C86000A4";
end if;
if first_state_sram_input_id = 1271 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1272 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1273 then
	sram_write <= x"44446000";
end if;
if first_state_sram_input_id = 1274 then
	sram_write <= x"C86000A0";
end if;
if first_state_sram_input_id = 1275 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1276 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1277 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1278 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1279 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 1280 then
	sram_write <= x"C860009C";
end if;
if first_state_sram_input_id = 1281 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1282 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1283 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1284 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1285 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1286 then
	sram_write <= x"48262000";
end if;
if first_state_sram_input_id = 1287 then
	sram_write <= x"44242000";
end if;
if first_state_sram_input_id = 1288 then
	sram_write <= x"8200147C";
end if;
if first_state_sram_input_id = 1289 then
	sram_write <= x"44262000";
end if;
if first_state_sram_input_id = 1290 then
	sram_write <= x"C84000B4";
end if;
if first_state_sram_input_id = 1291 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 1292 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 1293 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 1294 then
	sram_write <= x"44424000";
end if;
if first_state_sram_input_id = 1295 then
	sram_write <= x"C86000B0";
end if;
if first_state_sram_input_id = 1296 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1297 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1298 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1299 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1300 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1301 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 1302 then
	sram_write <= x"C86000AC";
end if;
if first_state_sram_input_id = 1303 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1304 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1305 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1306 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1307 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1308 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1309 then
	sram_write <= x"48262000";
end if;
if first_state_sram_input_id = 1310 then
	sram_write <= x"44242000";
end if;
if first_state_sram_input_id = 1311 then
	sram_write <= x"44202000";
end if;
if first_state_sram_input_id = 1312 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 1313 then
	sram_write <= x"C84000C0";
end if;
if first_state_sram_input_id = 1314 then
	sram_write <= x"C86000BC";
end if;
if first_state_sram_input_id = 1315 then
	sram_write <= x"C88000B8";
end if;
if first_state_sram_input_id = 1316 then
	sram_write <= x"8E2414B8";
end if;
if first_state_sram_input_id = 1317 then
	sram_write <= x"44224000";
end if;
if first_state_sram_input_id = 1318 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 1319 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1320 then
	sram_write <= x"03DC0008";
end if;
if first_state_sram_input_id = 1321 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1322 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1323 then
	sram_write <= x"8200084C";
end if;
if first_state_sram_input_id = 1324 then
	sram_write <= x"07DC0008";
end if;
if first_state_sram_input_id = 1325 then
	sram_write <= x"82001618";
end if;
if first_state_sram_input_id = 1326 then
	sram_write <= x"8E26156C";
end if;
if first_state_sram_input_id = 1327 then
	sram_write <= x"8E821510";
end if;
if first_state_sram_input_id = 1328 then
	sram_write <= x"C84000A8";
end if;
if first_state_sram_input_id = 1329 then
	sram_write <= x"C86000A4";
end if;
if first_state_sram_input_id = 1330 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1331 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1332 then
	sram_write <= x"44446000";
end if;
if first_state_sram_input_id = 1333 then
	sram_write <= x"C86000A0";
end if;
if first_state_sram_input_id = 1334 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1335 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1336 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1337 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1338 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 1339 then
	sram_write <= x"C860009C";
end if;
if first_state_sram_input_id = 1340 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1341 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1342 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1343 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1344 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1345 then
	sram_write <= x"48262000";
end if;
if first_state_sram_input_id = 1346 then
	sram_write <= x"44242000";
end if;
if first_state_sram_input_id = 1347 then
	sram_write <= x"82001568";
end if;
if first_state_sram_input_id = 1348 then
	sram_write <= x"44262000";
end if;
if first_state_sram_input_id = 1349 then
	sram_write <= x"C84000B4";
end if;
if first_state_sram_input_id = 1350 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 1351 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 1352 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 1353 then
	sram_write <= x"44424000";
end if;
if first_state_sram_input_id = 1354 then
	sram_write <= x"C86000B0";
end if;
if first_state_sram_input_id = 1355 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1356 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1357 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1358 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1359 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1360 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 1361 then
	sram_write <= x"C86000AC";
end if;
if first_state_sram_input_id = 1362 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1363 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1364 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1365 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1366 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1367 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1368 then
	sram_write <= x"48262000";
end if;
if first_state_sram_input_id = 1369 then
	sram_write <= x"44242000";
end if;
if first_state_sram_input_id = 1370 then
	sram_write <= x"82001618";
end if;
if first_state_sram_input_id = 1371 then
	sram_write <= x"8E8215C0";
end if;
if first_state_sram_input_id = 1372 then
	sram_write <= x"C84000A8";
end if;
if first_state_sram_input_id = 1373 then
	sram_write <= x"C86000A4";
end if;
if first_state_sram_input_id = 1374 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1375 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1376 then
	sram_write <= x"44446000";
end if;
if first_state_sram_input_id = 1377 then
	sram_write <= x"C86000A0";
end if;
if first_state_sram_input_id = 1378 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1379 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1380 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1381 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1382 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 1383 then
	sram_write <= x"C860009C";
end if;
if first_state_sram_input_id = 1384 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1385 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1386 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1387 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1388 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1389 then
	sram_write <= x"48262000";
end if;
if first_state_sram_input_id = 1390 then
	sram_write <= x"44242000";
end if;
if first_state_sram_input_id = 1391 then
	sram_write <= x"82001618";
end if;
if first_state_sram_input_id = 1392 then
	sram_write <= x"44262000";
end if;
if first_state_sram_input_id = 1393 then
	sram_write <= x"C84000B4";
end if;
if first_state_sram_input_id = 1394 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 1395 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 1396 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 1397 then
	sram_write <= x"44424000";
end if;
if first_state_sram_input_id = 1398 then
	sram_write <= x"C86000B0";
end if;
if first_state_sram_input_id = 1399 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1400 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1401 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1402 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1403 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1404 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 1405 then
	sram_write <= x"C86000AC";
end if;
if first_state_sram_input_id = 1406 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1407 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1408 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1409 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1410 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1411 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 1412 then
	sram_write <= x"48262000";
end if;
if first_state_sram_input_id = 1413 then
	sram_write <= x"44242000";
end if;
if first_state_sram_input_id = 1414 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 1415 then
	sram_write <= x"C8220000";
end if;
if first_state_sram_input_id = 1416 then
	sram_write <= x"48222000";
end if;
if first_state_sram_input_id = 1417 then
	sram_write <= x"C8420004";
end if;
if first_state_sram_input_id = 1418 then
	sram_write <= x"48444000";
end if;
if first_state_sram_input_id = 1419 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 1420 then
	sram_write <= x"C8420008";
end if;
if first_state_sram_input_id = 1421 then
	sram_write <= x"48444000";
end if;
if first_state_sram_input_id = 1422 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 1423 then
	sram_write <= x"C43C0000";
end if;
if first_state_sram_input_id = 1424 then
	sram_write <= x"C45C0004";
end if;
if first_state_sram_input_id = 1425 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1426 then
	sram_write <= x"03DC0010";
end if;
if first_state_sram_input_id = 1427 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1428 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1429 then
	sram_write <= x"8200083C";
end if;
if first_state_sram_input_id = 1430 then
	sram_write <= x"07DC0010";
end if;
if first_state_sram_input_id = 1431 then
	sram_write <= x"8A2016A4";
end if;
if first_state_sram_input_id = 1432 then
	sram_write <= x"C03C0004";
end if;
if first_state_sram_input_id = 1433 then
	sram_write <= x"82201688";
end if;
if first_state_sram_input_id = 1434 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1435 then
	sram_write <= x"03DC0010";
end if;
if first_state_sram_input_id = 1436 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1437 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1438 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 1439 then
	sram_write <= x"07DC0010";
end if;
if first_state_sram_input_id = 1440 then
	sram_write <= x"44202000";
end if;
if first_state_sram_input_id = 1441 then
	sram_write <= x"820016A0";
end if;
if first_state_sram_input_id = 1442 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1443 then
	sram_write <= x"03DC0010";
end if;
if first_state_sram_input_id = 1444 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1445 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1446 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 1447 then
	sram_write <= x"07DC0010";
end if;
if first_state_sram_input_id = 1448 then
	sram_write <= x"820016A8";
end if;
if first_state_sram_input_id = 1449 then
	sram_write <= x"C82000A8";
end if;
if first_state_sram_input_id = 1450 then
	sram_write <= x"C03C0000";
end if;
if first_state_sram_input_id = 1451 then
	sram_write <= x"C8420000";
end if;
if first_state_sram_input_id = 1452 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 1453 then
	sram_write <= x"CC420000";
end if;
if first_state_sram_input_id = 1454 then
	sram_write <= x"C8420004";
end if;
if first_state_sram_input_id = 1455 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 1456 then
	sram_write <= x"CC420004";
end if;
if first_state_sram_input_id = 1457 then
	sram_write <= x"C8420008";
end if;
if first_state_sram_input_id = 1458 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 1459 then
	sram_write <= x"CC220008";
end if;
if first_state_sram_input_id = 1460 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 1461 then
	sram_write <= x"022001B8";
end if;
if first_state_sram_input_id = 1462 then
	sram_write <= x"C43C0000";
end if;
if first_state_sram_input_id = 1463 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1464 then
	sram_write <= x"03DC000C";
end if;
if first_state_sram_input_id = 1465 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1466 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1467 then
	sram_write <= x"820007C0";
end if;
if first_state_sram_input_id = 1468 then
	sram_write <= x"07DC000C";
end if;
if first_state_sram_input_id = 1469 then
	sram_write <= x"C03C0000";
end if;
if first_state_sram_input_id = 1470 then
	sram_write <= x"CC220000";
end if;
if first_state_sram_input_id = 1471 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1472 then
	sram_write <= x"03DC000C";
end if;
if first_state_sram_input_id = 1473 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1474 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1475 then
	sram_write <= x"820007C0";
end if;
if first_state_sram_input_id = 1476 then
	sram_write <= x"07DC000C";
end if;
if first_state_sram_input_id = 1477 then
	sram_write <= x"C03C0000";
end if;
if first_state_sram_input_id = 1478 then
	sram_write <= x"CC220004";
end if;
if first_state_sram_input_id = 1479 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1480 then
	sram_write <= x"03DC000C";
end if;
if first_state_sram_input_id = 1481 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1482 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1483 then
	sram_write <= x"820007C0";
end if;
if first_state_sram_input_id = 1484 then
	sram_write <= x"07DC000C";
end if;
if first_state_sram_input_id = 1485 then
	sram_write <= x"C03C0000";
end if;
if first_state_sram_input_id = 1486 then
	sram_write <= x"CC220008";
end if;
if first_state_sram_input_id = 1487 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1488 then
	sram_write <= x"03DC000C";
end if;
if first_state_sram_input_id = 1489 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1490 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1491 then
	sram_write <= x"820007C0";
end if;
if first_state_sram_input_id = 1492 then
	sram_write <= x"07DC000C";
end if;
if first_state_sram_input_id = 1493 then
	sram_write <= x"C840008C";
end if;
if first_state_sram_input_id = 1494 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 1495 then
	sram_write <= x"C8600098";
end if;
if first_state_sram_input_id = 1496 then
	sram_write <= x"CC5C0008";
end if;
if first_state_sram_input_id = 1497 then
	sram_write <= x"CC7C0010";
end if;
if first_state_sram_input_id = 1498 then
	sram_write <= x"CC3C0018";
end if;
if first_state_sram_input_id = 1499 then
	sram_write <= x"8E261794";
end if;
if first_state_sram_input_id = 1500 then
	sram_write <= x"44826000";
end if;
if first_state_sram_input_id = 1501 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1502 then
	sram_write <= x"40208000";
end if;
if first_state_sram_input_id = 1503 then
	sram_write <= x"03DC0028";
end if;
if first_state_sram_input_id = 1504 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1505 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1506 then
	sram_write <= x"82001270";
end if;
if first_state_sram_input_id = 1507 then
	sram_write <= x"07DC0028";
end if;
if first_state_sram_input_id = 1508 then
	sram_write <= x"82001800";
end if;
if first_state_sram_input_id = 1509 then
	sram_write <= x"8E0217E4";
end if;
if first_state_sram_input_id = 1510 then
	sram_write <= x"C8800090";
end if;
if first_state_sram_input_id = 1511 then
	sram_write <= x"8E8217C4";
end if;
if first_state_sram_input_id = 1512 then
	sram_write <= x"40826000";
end if;
if first_state_sram_input_id = 1513 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1514 then
	sram_write <= x"40208000";
end if;
if first_state_sram_input_id = 1515 then
	sram_write <= x"03DC0028";
end if;
if first_state_sram_input_id = 1516 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1517 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1518 then
	sram_write <= x"82001270";
end if;
if first_state_sram_input_id = 1519 then
	sram_write <= x"07DC0028";
end if;
if first_state_sram_input_id = 1520 then
	sram_write <= x"820017E0";
end if;
if first_state_sram_input_id = 1521 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 1522 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1523 then
	sram_write <= x"03DC0028";
end if;
if first_state_sram_input_id = 1524 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1525 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1526 then
	sram_write <= x"82000B88";
end if;
if first_state_sram_input_id = 1527 then
	sram_write <= x"07DC0028";
end if;
if first_state_sram_input_id = 1528 then
	sram_write <= x"82001800";
end if;
if first_state_sram_input_id = 1529 then
	sram_write <= x"0220FFFF";
end if;
if first_state_sram_input_id = 1530 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1531 then
	sram_write <= x"03DC0028";
end if;
if first_state_sram_input_id = 1532 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1533 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1534 then
	sram_write <= x"82000B88";
end if;
if first_state_sram_input_id = 1535 then
	sram_write <= x"07DC0028";
end if;
if first_state_sram_input_id = 1536 then
	sram_write <= x"C85C0010";
end if;
if first_state_sram_input_id = 1537 then
	sram_write <= x"C87C0018";
end if;
if first_state_sram_input_id = 1538 then
	sram_write <= x"CC3C0020";
end if;
if first_state_sram_input_id = 1539 then
	sram_write <= x"8E641834";
end if;
if first_state_sram_input_id = 1540 then
	sram_write <= x"44664000";
end if;
if first_state_sram_input_id = 1541 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1542 then
	sram_write <= x"40206000";
end if;
if first_state_sram_input_id = 1543 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 1544 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1545 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1546 then
	sram_write <= x"82000EC4";
end if;
if first_state_sram_input_id = 1547 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 1548 then
	sram_write <= x"820018A8";
end if;
if first_state_sram_input_id = 1549 then
	sram_write <= x"8E061888";
end if;
if first_state_sram_input_id = 1550 then
	sram_write <= x"C8800090";
end if;
if first_state_sram_input_id = 1551 then
	sram_write <= x"8E861864";
end if;
if first_state_sram_input_id = 1552 then
	sram_write <= x"40664000";
end if;
if first_state_sram_input_id = 1553 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1554 then
	sram_write <= x"40206000";
end if;
if first_state_sram_input_id = 1555 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 1556 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1557 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1558 then
	sram_write <= x"82000EC4";
end if;
if first_state_sram_input_id = 1559 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 1560 then
	sram_write <= x"82001884";
end if;
if first_state_sram_input_id = 1561 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 1562 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1563 then
	sram_write <= x"40206000";
end if;
if first_state_sram_input_id = 1564 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 1565 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1566 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1567 then
	sram_write <= x"8200084C";
end if;
if first_state_sram_input_id = 1568 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 1569 then
	sram_write <= x"820018A8";
end if;
if first_state_sram_input_id = 1570 then
	sram_write <= x"0220FFFF";
end if;
if first_state_sram_input_id = 1571 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1572 then
	sram_write <= x"40206000";
end if;
if first_state_sram_input_id = 1573 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 1574 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1575 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1576 then
	sram_write <= x"8200084C";
end if;
if first_state_sram_input_id = 1577 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 1578 then
	sram_write <= x"CC3C0028";
end if;
if first_state_sram_input_id = 1579 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1580 then
	sram_write <= x"03DC0038";
end if;
if first_state_sram_input_id = 1581 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1582 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1583 then
	sram_write <= x"820007C0";
end if;
if first_state_sram_input_id = 1584 then
	sram_write <= x"07DC0038";
end if;
if first_state_sram_input_id = 1585 then
	sram_write <= x"C85C0008";
end if;
if first_state_sram_input_id = 1586 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 1587 then
	sram_write <= x"C85C0010";
end if;
if first_state_sram_input_id = 1588 then
	sram_write <= x"CC3C0030";
end if;
if first_state_sram_input_id = 1589 then
	sram_write <= x"8E2418FC";
end if;
if first_state_sram_input_id = 1590 then
	sram_write <= x"44624000";
end if;
if first_state_sram_input_id = 1591 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1592 then
	sram_write <= x"40206000";
end if;
if first_state_sram_input_id = 1593 then
	sram_write <= x"03DC0040";
end if;
if first_state_sram_input_id = 1594 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1595 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1596 then
	sram_write <= x"82001270";
end if;
if first_state_sram_input_id = 1597 then
	sram_write <= x"07DC0040";
end if;
if first_state_sram_input_id = 1598 then
	sram_write <= x"82001968";
end if;
if first_state_sram_input_id = 1599 then
	sram_write <= x"8E02194C";
end if;
if first_state_sram_input_id = 1600 then
	sram_write <= x"C8600090";
end if;
if first_state_sram_input_id = 1601 then
	sram_write <= x"8E62192C";
end if;
if first_state_sram_input_id = 1602 then
	sram_write <= x"40624000";
end if;
if first_state_sram_input_id = 1603 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1604 then
	sram_write <= x"40206000";
end if;
if first_state_sram_input_id = 1605 then
	sram_write <= x"03DC0040";
end if;
if first_state_sram_input_id = 1606 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1607 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1608 then
	sram_write <= x"82001270";
end if;
if first_state_sram_input_id = 1609 then
	sram_write <= x"07DC0040";
end if;
if first_state_sram_input_id = 1610 then
	sram_write <= x"82001948";
end if;
if first_state_sram_input_id = 1611 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 1612 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1613 then
	sram_write <= x"03DC0040";
end if;
if first_state_sram_input_id = 1614 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1615 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1616 then
	sram_write <= x"82000B88";
end if;
if first_state_sram_input_id = 1617 then
	sram_write <= x"07DC0040";
end if;
if first_state_sram_input_id = 1618 then
	sram_write <= x"82001968";
end if;
if first_state_sram_input_id = 1619 then
	sram_write <= x"0220FFFF";
end if;
if first_state_sram_input_id = 1620 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1621 then
	sram_write <= x"03DC0040";
end if;
if first_state_sram_input_id = 1622 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1623 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1624 then
	sram_write <= x"82000B88";
end if;
if first_state_sram_input_id = 1625 then
	sram_write <= x"07DC0040";
end if;
if first_state_sram_input_id = 1626 then
	sram_write <= x"C85C0010";
end if;
if first_state_sram_input_id = 1627 then
	sram_write <= x"C87C0030";
end if;
if first_state_sram_input_id = 1628 then
	sram_write <= x"CC3C0038";
end if;
if first_state_sram_input_id = 1629 then
	sram_write <= x"8E64199C";
end if;
if first_state_sram_input_id = 1630 then
	sram_write <= x"44464000";
end if;
if first_state_sram_input_id = 1631 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1632 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 1633 then
	sram_write <= x"03DC0048";
end if;
if first_state_sram_input_id = 1634 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1635 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1636 then
	sram_write <= x"82000EC4";
end if;
if first_state_sram_input_id = 1637 then
	sram_write <= x"07DC0048";
end if;
if first_state_sram_input_id = 1638 then
	sram_write <= x"82001A10";
end if;
if first_state_sram_input_id = 1639 then
	sram_write <= x"8E0619F0";
end if;
if first_state_sram_input_id = 1640 then
	sram_write <= x"C8800090";
end if;
if first_state_sram_input_id = 1641 then
	sram_write <= x"8E8619CC";
end if;
if first_state_sram_input_id = 1642 then
	sram_write <= x"40464000";
end if;
if first_state_sram_input_id = 1643 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1644 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 1645 then
	sram_write <= x"03DC0048";
end if;
if first_state_sram_input_id = 1646 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1647 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1648 then
	sram_write <= x"82000EC4";
end if;
if first_state_sram_input_id = 1649 then
	sram_write <= x"07DC0048";
end if;
if first_state_sram_input_id = 1650 then
	sram_write <= x"820019EC";
end if;
if first_state_sram_input_id = 1651 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 1652 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1653 then
	sram_write <= x"40206000";
end if;
if first_state_sram_input_id = 1654 then
	sram_write <= x"03DC0048";
end if;
if first_state_sram_input_id = 1655 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1656 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1657 then
	sram_write <= x"8200084C";
end if;
if first_state_sram_input_id = 1658 then
	sram_write <= x"07DC0048";
end if;
if first_state_sram_input_id = 1659 then
	sram_write <= x"82001A10";
end if;
if first_state_sram_input_id = 1660 then
	sram_write <= x"0220FFFF";
end if;
if first_state_sram_input_id = 1661 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1662 then
	sram_write <= x"40206000";
end if;
if first_state_sram_input_id = 1663 then
	sram_write <= x"03DC0048";
end if;
if first_state_sram_input_id = 1664 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1665 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1666 then
	sram_write <= x"8200084C";
end if;
if first_state_sram_input_id = 1667 then
	sram_write <= x"07DC0048";
end if;
if first_state_sram_input_id = 1668 then
	sram_write <= x"0220033C";
end if;
if first_state_sram_input_id = 1669 then
	sram_write <= x"C85C0020";
end if;
if first_state_sram_input_id = 1670 then
	sram_write <= x"48642000";
end if;
if first_state_sram_input_id = 1671 then
	sram_write <= x"C8800088";
end if;
if first_state_sram_input_id = 1672 then
	sram_write <= x"48668000";
end if;
if first_state_sram_input_id = 1673 then
	sram_write <= x"CC620000";
end if;
if first_state_sram_input_id = 1674 then
	sram_write <= x"C8600084";
end if;
if first_state_sram_input_id = 1675 then
	sram_write <= x"C8BC0028";
end if;
if first_state_sram_input_id = 1676 then
	sram_write <= x"486A6000";
end if;
if first_state_sram_input_id = 1677 then
	sram_write <= x"CC620004";
end if;
if first_state_sram_input_id = 1678 then
	sram_write <= x"C87C0038";
end if;
if first_state_sram_input_id = 1679 then
	sram_write <= x"48C46000";
end if;
if first_state_sram_input_id = 1680 then
	sram_write <= x"488C8000";
end if;
if first_state_sram_input_id = 1681 then
	sram_write <= x"CC820008";
end if;
if first_state_sram_input_id = 1682 then
	sram_write <= x"02400324";
end if;
if first_state_sram_input_id = 1683 then
	sram_write <= x"CC640000";
end if;
if first_state_sram_input_id = 1684 then
	sram_write <= x"CC040004";
end if;
if first_state_sram_input_id = 1685 then
	sram_write <= x"44802000";
end if;
if first_state_sram_input_id = 1686 then
	sram_write <= x"CC840008";
end if;
if first_state_sram_input_id = 1687 then
	sram_write <= x"02400330";
end if;
if first_state_sram_input_id = 1688 then
	sram_write <= x"4480A000";
end if;
if first_state_sram_input_id = 1689 then
	sram_write <= x"48282000";
end if;
if first_state_sram_input_id = 1690 then
	sram_write <= x"CC240000";
end if;
if first_state_sram_input_id = 1691 then
	sram_write <= x"44204000";
end if;
if first_state_sram_input_id = 1692 then
	sram_write <= x"CC240004";
end if;
if first_state_sram_input_id = 1693 then
	sram_write <= x"48286000";
end if;
if first_state_sram_input_id = 1694 then
	sram_write <= x"CC240008";
end if;
if first_state_sram_input_id = 1695 then
	sram_write <= x"024001C4";
end if;
if first_state_sram_input_id = 1696 then
	sram_write <= x"C07C0000";
end if;
if first_state_sram_input_id = 1697 then
	sram_write <= x"C8260000";
end if;
if first_state_sram_input_id = 1698 then
	sram_write <= x"C8420000";
end if;
if first_state_sram_input_id = 1699 then
	sram_write <= x"44224000";
end if;
if first_state_sram_input_id = 1700 then
	sram_write <= x"CC240000";
end if;
if first_state_sram_input_id = 1701 then
	sram_write <= x"C8260004";
end if;
if first_state_sram_input_id = 1702 then
	sram_write <= x"C8420004";
end if;
if first_state_sram_input_id = 1703 then
	sram_write <= x"44224000";
end if;
if first_state_sram_input_id = 1704 then
	sram_write <= x"CC240004";
end if;
if first_state_sram_input_id = 1705 then
	sram_write <= x"C8260008";
end if;
if first_state_sram_input_id = 1706 then
	sram_write <= x"C8420008";
end if;
if first_state_sram_input_id = 1707 then
	sram_write <= x"44224000";
end if;
if first_state_sram_input_id = 1708 then
	sram_write <= x"CC240008";
end if;
if first_state_sram_input_id = 1709 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 1710 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1711 then
	sram_write <= x"03DC0008";
end if;
if first_state_sram_input_id = 1712 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1713 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1714 then
	sram_write <= x"82000794";
end if;
if first_state_sram_input_id = 1715 then
	sram_write <= x"07DC0008";
end if;
if first_state_sram_input_id = 1716 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1717 then
	sram_write <= x"03DC0008";
end if;
if first_state_sram_input_id = 1718 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1719 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1720 then
	sram_write <= x"820007C0";
end if;
if first_state_sram_input_id = 1721 then
	sram_write <= x"07DC0008";
end if;
if first_state_sram_input_id = 1722 then
	sram_write <= x"C840008C";
end if;
if first_state_sram_input_id = 1723 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 1724 then
	sram_write <= x"C8600098";
end if;
if first_state_sram_input_id = 1725 then
	sram_write <= x"CC7C0000";
end if;
if first_state_sram_input_id = 1726 then
	sram_write <= x"CC3C0008";
end if;
if first_state_sram_input_id = 1727 then
	sram_write <= x"CC5C0010";
end if;
if first_state_sram_input_id = 1728 then
	sram_write <= x"8E261B28";
end if;
if first_state_sram_input_id = 1729 then
	sram_write <= x"44826000";
end if;
if first_state_sram_input_id = 1730 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1731 then
	sram_write <= x"40208000";
end if;
if first_state_sram_input_id = 1732 then
	sram_write <= x"03DC0020";
end if;
if first_state_sram_input_id = 1733 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1734 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1735 then
	sram_write <= x"82000EC4";
end if;
if first_state_sram_input_id = 1736 then
	sram_write <= x"07DC0020";
end if;
if first_state_sram_input_id = 1737 then
	sram_write <= x"82001B94";
end if;
if first_state_sram_input_id = 1738 then
	sram_write <= x"8E021B78";
end if;
if first_state_sram_input_id = 1739 then
	sram_write <= x"C8800090";
end if;
if first_state_sram_input_id = 1740 then
	sram_write <= x"8E821B58";
end if;
if first_state_sram_input_id = 1741 then
	sram_write <= x"40826000";
end if;
if first_state_sram_input_id = 1742 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1743 then
	sram_write <= x"40208000";
end if;
if first_state_sram_input_id = 1744 then
	sram_write <= x"03DC0020";
end if;
if first_state_sram_input_id = 1745 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1746 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1747 then
	sram_write <= x"82000EC4";
end if;
if first_state_sram_input_id = 1748 then
	sram_write <= x"07DC0020";
end if;
if first_state_sram_input_id = 1749 then
	sram_write <= x"82001B74";
end if;
if first_state_sram_input_id = 1750 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 1751 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1752 then
	sram_write <= x"03DC0020";
end if;
if first_state_sram_input_id = 1753 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1754 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1755 then
	sram_write <= x"8200084C";
end if;
if first_state_sram_input_id = 1756 then
	sram_write <= x"07DC0020";
end if;
if first_state_sram_input_id = 1757 then
	sram_write <= x"82001B94";
end if;
if first_state_sram_input_id = 1758 then
	sram_write <= x"0220FFFF";
end if;
if first_state_sram_input_id = 1759 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1760 then
	sram_write <= x"03DC0020";
end if;
if first_state_sram_input_id = 1761 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1762 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1763 then
	sram_write <= x"8200084C";
end if;
if first_state_sram_input_id = 1764 then
	sram_write <= x"07DC0020";
end if;
if first_state_sram_input_id = 1765 then
	sram_write <= x"022001D0";
end if;
if first_state_sram_input_id = 1766 then
	sram_write <= x"44202000";
end if;
if first_state_sram_input_id = 1767 then
	sram_write <= x"CC220004";
end if;
if first_state_sram_input_id = 1768 then
	sram_write <= x"C43C0018";
end if;
if first_state_sram_input_id = 1769 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1770 then
	sram_write <= x"03DC0024";
end if;
if first_state_sram_input_id = 1771 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1772 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1773 then
	sram_write <= x"820007C0";
end if;
if first_state_sram_input_id = 1774 then
	sram_write <= x"07DC0024";
end if;
if first_state_sram_input_id = 1775 then
	sram_write <= x"C85C0010";
end if;
if first_state_sram_input_id = 1776 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 1777 then
	sram_write <= x"C85C0000";
end if;
if first_state_sram_input_id = 1778 then
	sram_write <= x"C87C0008";
end if;
if first_state_sram_input_id = 1779 then
	sram_write <= x"CC3C0020";
end if;
if first_state_sram_input_id = 1780 then
	sram_write <= x"8E641BF8";
end if;
if first_state_sram_input_id = 1781 then
	sram_write <= x"44664000";
end if;
if first_state_sram_input_id = 1782 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1783 then
	sram_write <= x"40206000";
end if;
if first_state_sram_input_id = 1784 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 1785 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1786 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1787 then
	sram_write <= x"82001270";
end if;
if first_state_sram_input_id = 1788 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 1789 then
	sram_write <= x"82001C6C";
end if;
if first_state_sram_input_id = 1790 then
	sram_write <= x"8E061C4C";
end if;
if first_state_sram_input_id = 1791 then
	sram_write <= x"C8800090";
end if;
if first_state_sram_input_id = 1792 then
	sram_write <= x"8E861C28";
end if;
if first_state_sram_input_id = 1793 then
	sram_write <= x"40664000";
end if;
if first_state_sram_input_id = 1794 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1795 then
	sram_write <= x"40206000";
end if;
if first_state_sram_input_id = 1796 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 1797 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1798 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1799 then
	sram_write <= x"82001270";
end if;
if first_state_sram_input_id = 1800 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 1801 then
	sram_write <= x"82001C48";
end if;
if first_state_sram_input_id = 1802 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 1803 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1804 then
	sram_write <= x"40206000";
end if;
if first_state_sram_input_id = 1805 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 1806 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1807 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1808 then
	sram_write <= x"82000B88";
end if;
if first_state_sram_input_id = 1809 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 1810 then
	sram_write <= x"82001C6C";
end if;
if first_state_sram_input_id = 1811 then
	sram_write <= x"0220FFFF";
end if;
if first_state_sram_input_id = 1812 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1813 then
	sram_write <= x"40206000";
end if;
if first_state_sram_input_id = 1814 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 1815 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1816 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1817 then
	sram_write <= x"82000B88";
end if;
if first_state_sram_input_id = 1818 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 1819 then
	sram_write <= x"C85C0000";
end if;
if first_state_sram_input_id = 1820 then
	sram_write <= x"C87C0020";
end if;
if first_state_sram_input_id = 1821 then
	sram_write <= x"CC3C0028";
end if;
if first_state_sram_input_id = 1822 then
	sram_write <= x"8E641CA0";
end if;
if first_state_sram_input_id = 1823 then
	sram_write <= x"44864000";
end if;
if first_state_sram_input_id = 1824 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1825 then
	sram_write <= x"40208000";
end if;
if first_state_sram_input_id = 1826 then
	sram_write <= x"03DC0038";
end if;
if first_state_sram_input_id = 1827 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1828 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1829 then
	sram_write <= x"82000EC4";
end if;
if first_state_sram_input_id = 1830 then
	sram_write <= x"07DC0038";
end if;
if first_state_sram_input_id = 1831 then
	sram_write <= x"82001D14";
end if;
if first_state_sram_input_id = 1832 then
	sram_write <= x"8E061CF4";
end if;
if first_state_sram_input_id = 1833 then
	sram_write <= x"C8800090";
end if;
if first_state_sram_input_id = 1834 then
	sram_write <= x"8E861CD0";
end if;
if first_state_sram_input_id = 1835 then
	sram_write <= x"40864000";
end if;
if first_state_sram_input_id = 1836 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1837 then
	sram_write <= x"40208000";
end if;
if first_state_sram_input_id = 1838 then
	sram_write <= x"03DC0038";
end if;
if first_state_sram_input_id = 1839 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1840 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1841 then
	sram_write <= x"82000EC4";
end if;
if first_state_sram_input_id = 1842 then
	sram_write <= x"07DC0038";
end if;
if first_state_sram_input_id = 1843 then
	sram_write <= x"82001CF0";
end if;
if first_state_sram_input_id = 1844 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 1845 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1846 then
	sram_write <= x"40206000";
end if;
if first_state_sram_input_id = 1847 then
	sram_write <= x"03DC0038";
end if;
if first_state_sram_input_id = 1848 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1849 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1850 then
	sram_write <= x"8200084C";
end if;
if first_state_sram_input_id = 1851 then
	sram_write <= x"07DC0038";
end if;
if first_state_sram_input_id = 1852 then
	sram_write <= x"82001D14";
end if;
if first_state_sram_input_id = 1853 then
	sram_write <= x"0220FFFF";
end if;
if first_state_sram_input_id = 1854 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1855 then
	sram_write <= x"40206000";
end if;
if first_state_sram_input_id = 1856 then
	sram_write <= x"03DC0038";
end if;
if first_state_sram_input_id = 1857 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1858 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1859 then
	sram_write <= x"8200084C";
end if;
if first_state_sram_input_id = 1860 then
	sram_write <= x"07DC0038";
end if;
if first_state_sram_input_id = 1861 then
	sram_write <= x"C85C0028";
end if;
if first_state_sram_input_id = 1862 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 1863 then
	sram_write <= x"C03C0018";
end if;
if first_state_sram_input_id = 1864 then
	sram_write <= x"CC220000";
end if;
if first_state_sram_input_id = 1865 then
	sram_write <= x"C83C0000";
end if;
if first_state_sram_input_id = 1866 then
	sram_write <= x"C87C0020";
end if;
if first_state_sram_input_id = 1867 then
	sram_write <= x"8E621D50";
end if;
if first_state_sram_input_id = 1868 then
	sram_write <= x"44262000";
end if;
if first_state_sram_input_id = 1869 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1870 then
	sram_write <= x"03DC0038";
end if;
if first_state_sram_input_id = 1871 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1872 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1873 then
	sram_write <= x"82001270";
end if;
if first_state_sram_input_id = 1874 then
	sram_write <= x"07DC0038";
end if;
if first_state_sram_input_id = 1875 then
	sram_write <= x"82001DC8";
end if;
if first_state_sram_input_id = 1876 then
	sram_write <= x"8E061DA4";
end if;
if first_state_sram_input_id = 1877 then
	sram_write <= x"C8800090";
end if;
if first_state_sram_input_id = 1878 then
	sram_write <= x"8E861D7C";
end if;
if first_state_sram_input_id = 1879 then
	sram_write <= x"40262000";
end if;
if first_state_sram_input_id = 1880 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1881 then
	sram_write <= x"03DC0038";
end if;
if first_state_sram_input_id = 1882 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1883 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1884 then
	sram_write <= x"82001270";
end if;
if first_state_sram_input_id = 1885 then
	sram_write <= x"07DC0038";
end if;
if first_state_sram_input_id = 1886 then
	sram_write <= x"82001DA0";
end if;
if first_state_sram_input_id = 1887 then
	sram_write <= x"02400001";
end if;
if first_state_sram_input_id = 1888 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1889 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 1890 then
	sram_write <= x"40206000";
end if;
if first_state_sram_input_id = 1891 then
	sram_write <= x"03DC0038";
end if;
if first_state_sram_input_id = 1892 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1893 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1894 then
	sram_write <= x"82000B88";
end if;
if first_state_sram_input_id = 1895 then
	sram_write <= x"07DC0038";
end if;
if first_state_sram_input_id = 1896 then
	sram_write <= x"82001DC8";
end if;
if first_state_sram_input_id = 1897 then
	sram_write <= x"0240FFFF";
end if;
if first_state_sram_input_id = 1898 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1899 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 1900 then
	sram_write <= x"40206000";
end if;
if first_state_sram_input_id = 1901 then
	sram_write <= x"03DC0038";
end if;
if first_state_sram_input_id = 1902 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1903 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1904 then
	sram_write <= x"82000B88";
end if;
if first_state_sram_input_id = 1905 then
	sram_write <= x"07DC0038";
end if;
if first_state_sram_input_id = 1906 then
	sram_write <= x"C85C0028";
end if;
if first_state_sram_input_id = 1907 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 1908 then
	sram_write <= x"C03C0018";
end if;
if first_state_sram_input_id = 1909 then
	sram_write <= x"CC220008";
end if;
if first_state_sram_input_id = 1910 then
	sram_write <= x"022001DC";
end if;
if first_state_sram_input_id = 1911 then
	sram_write <= x"C43C0030";
end if;
if first_state_sram_input_id = 1912 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1913 then
	sram_write <= x"03DC003C";
end if;
if first_state_sram_input_id = 1914 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1915 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1916 then
	sram_write <= x"820007C0";
end if;
if first_state_sram_input_id = 1917 then
	sram_write <= x"07DC003C";
end if;
if first_state_sram_input_id = 1918 then
	sram_write <= x"C03C0030";
end if;
if first_state_sram_input_id = 1919 then
	sram_write <= x"CC220000";
end if;
if first_state_sram_input_id = 1920 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 1921 then
	sram_write <= x"C8240000";
end if;
if first_state_sram_input_id = 1922 then
	sram_write <= x"C8400098";
end if;
if first_state_sram_input_id = 1923 then
	sram_write <= x"C43C0000";
end if;
if first_state_sram_input_id = 1924 then
	sram_write <= x"CC5C0008";
end if;
if first_state_sram_input_id = 1925 then
	sram_write <= x"C45C0010";
end if;
if first_state_sram_input_id = 1926 then
	sram_write <= x"8E241E3C";
end if;
if first_state_sram_input_id = 1927 then
	sram_write <= x"44224000";
end if;
if first_state_sram_input_id = 1928 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1929 then
	sram_write <= x"03DC001C";
end if;
if first_state_sram_input_id = 1930 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1931 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1932 then
	sram_write <= x"82001270";
end if;
if first_state_sram_input_id = 1933 then
	sram_write <= x"07DC001C";
end if;
if first_state_sram_input_id = 1934 then
	sram_write <= x"82001EAC";
end if;
if first_state_sram_input_id = 1935 then
	sram_write <= x"8E021E8C";
end if;
if first_state_sram_input_id = 1936 then
	sram_write <= x"C8600090";
end if;
if first_state_sram_input_id = 1937 then
	sram_write <= x"8E621E68";
end if;
if first_state_sram_input_id = 1938 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 1939 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1940 then
	sram_write <= x"03DC001C";
end if;
if first_state_sram_input_id = 1941 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1942 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1943 then
	sram_write <= x"82001270";
end if;
if first_state_sram_input_id = 1944 then
	sram_write <= x"07DC001C";
end if;
if first_state_sram_input_id = 1945 then
	sram_write <= x"82001E88";
end if;
if first_state_sram_input_id = 1946 then
	sram_write <= x"02600001";
end if;
if first_state_sram_input_id = 1947 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1948 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 1949 then
	sram_write <= x"03DC001C";
end if;
if first_state_sram_input_id = 1950 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1951 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1952 then
	sram_write <= x"82000B88";
end if;
if first_state_sram_input_id = 1953 then
	sram_write <= x"07DC001C";
end if;
if first_state_sram_input_id = 1954 then
	sram_write <= x"82001EAC";
end if;
if first_state_sram_input_id = 1955 then
	sram_write <= x"0260FFFF";
end if;
if first_state_sram_input_id = 1956 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1957 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 1958 then
	sram_write <= x"03DC001C";
end if;
if first_state_sram_input_id = 1959 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1960 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1961 then
	sram_write <= x"82000B88";
end if;
if first_state_sram_input_id = 1962 then
	sram_write <= x"07DC001C";
end if;
if first_state_sram_input_id = 1963 then
	sram_write <= x"C03C0010";
end if;
if first_state_sram_input_id = 1964 then
	sram_write <= x"C8420000";
end if;
if first_state_sram_input_id = 1965 then
	sram_write <= x"C87C0008";
end if;
if first_state_sram_input_id = 1966 then
	sram_write <= x"CC3C0018";
end if;
if first_state_sram_input_id = 1967 then
	sram_write <= x"8E461EE4";
end if;
if first_state_sram_input_id = 1968 then
	sram_write <= x"44446000";
end if;
if first_state_sram_input_id = 1969 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1970 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 1971 then
	sram_write <= x"03DC0028";
end if;
if first_state_sram_input_id = 1972 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1973 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1974 then
	sram_write <= x"82000EC4";
end if;
if first_state_sram_input_id = 1975 then
	sram_write <= x"07DC0028";
end if;
if first_state_sram_input_id = 1976 then
	sram_write <= x"82001F60";
end if;
if first_state_sram_input_id = 1977 then
	sram_write <= x"8E041F3C";
end if;
if first_state_sram_input_id = 1978 then
	sram_write <= x"C8800090";
end if;
if first_state_sram_input_id = 1979 then
	sram_write <= x"8E841F14";
end if;
if first_state_sram_input_id = 1980 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 1981 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1982 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 1983 then
	sram_write <= x"03DC0028";
end if;
if first_state_sram_input_id = 1984 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1985 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1986 then
	sram_write <= x"82000EC4";
end if;
if first_state_sram_input_id = 1987 then
	sram_write <= x"07DC0028";
end if;
if first_state_sram_input_id = 1988 then
	sram_write <= x"82001F38";
end if;
if first_state_sram_input_id = 1989 then
	sram_write <= x"02400001";
end if;
if first_state_sram_input_id = 1990 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 1991 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 1992 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 1993 then
	sram_write <= x"03DC0028";
end if;
if first_state_sram_input_id = 1994 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 1995 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 1996 then
	sram_write <= x"8200084C";
end if;
if first_state_sram_input_id = 1997 then
	sram_write <= x"07DC0028";
end if;
if first_state_sram_input_id = 1998 then
	sram_write <= x"82001F60";
end if;
if first_state_sram_input_id = 1999 then
	sram_write <= x"0240FFFF";
end if;
if first_state_sram_input_id = 2000 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2001 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 2002 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 2003 then
	sram_write <= x"03DC0028";
end if;
if first_state_sram_input_id = 2004 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2005 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2006 then
	sram_write <= x"8200084C";
end if;
if first_state_sram_input_id = 2007 then
	sram_write <= x"07DC0028";
end if;
if first_state_sram_input_id = 2008 then
	sram_write <= x"C03C0010";
end if;
if first_state_sram_input_id = 2009 then
	sram_write <= x"C8420004";
end if;
if first_state_sram_input_id = 2010 then
	sram_write <= x"C87C0008";
end if;
if first_state_sram_input_id = 2011 then
	sram_write <= x"CC3C0020";
end if;
if first_state_sram_input_id = 2012 then
	sram_write <= x"8E461F98";
end if;
if first_state_sram_input_id = 2013 then
	sram_write <= x"44446000";
end if;
if first_state_sram_input_id = 2014 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2015 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 2016 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 2017 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2018 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2019 then
	sram_write <= x"82001270";
end if;
if first_state_sram_input_id = 2020 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 2021 then
	sram_write <= x"82002014";
end if;
if first_state_sram_input_id = 2022 then
	sram_write <= x"8E041FF0";
end if;
if first_state_sram_input_id = 2023 then
	sram_write <= x"C8800090";
end if;
if first_state_sram_input_id = 2024 then
	sram_write <= x"8E841FC8";
end if;
if first_state_sram_input_id = 2025 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 2026 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2027 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 2028 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 2029 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2030 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2031 then
	sram_write <= x"82001270";
end if;
if first_state_sram_input_id = 2032 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 2033 then
	sram_write <= x"82001FEC";
end if;
if first_state_sram_input_id = 2034 then
	sram_write <= x"02400001";
end if;
if first_state_sram_input_id = 2035 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2036 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 2037 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 2038 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 2039 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2040 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2041 then
	sram_write <= x"82000B88";
end if;
if first_state_sram_input_id = 2042 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 2043 then
	sram_write <= x"82002014";
end if;
if first_state_sram_input_id = 2044 then
	sram_write <= x"0240FFFF";
end if;
if first_state_sram_input_id = 2045 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2046 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 2047 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 2048 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 2049 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2050 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2051 then
	sram_write <= x"82000B88";
end if;
if first_state_sram_input_id = 2052 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 2053 then
	sram_write <= x"C03C0010";
end if;
if first_state_sram_input_id = 2054 then
	sram_write <= x"C8420004";
end if;
if first_state_sram_input_id = 2055 then
	sram_write <= x"C87C0008";
end if;
if first_state_sram_input_id = 2056 then
	sram_write <= x"CC3C0028";
end if;
if first_state_sram_input_id = 2057 then
	sram_write <= x"8E46204C";
end if;
if first_state_sram_input_id = 2058 then
	sram_write <= x"44446000";
end if;
if first_state_sram_input_id = 2059 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2060 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 2061 then
	sram_write <= x"03DC0038";
end if;
if first_state_sram_input_id = 2062 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2063 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2064 then
	sram_write <= x"82000EC4";
end if;
if first_state_sram_input_id = 2065 then
	sram_write <= x"07DC0038";
end if;
if first_state_sram_input_id = 2066 then
	sram_write <= x"820020C8";
end if;
if first_state_sram_input_id = 2067 then
	sram_write <= x"8E0420A4";
end if;
if first_state_sram_input_id = 2068 then
	sram_write <= x"C8800090";
end if;
if first_state_sram_input_id = 2069 then
	sram_write <= x"8E84207C";
end if;
if first_state_sram_input_id = 2070 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 2071 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2072 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 2073 then
	sram_write <= x"03DC0038";
end if;
if first_state_sram_input_id = 2074 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2075 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2076 then
	sram_write <= x"82000EC4";
end if;
if first_state_sram_input_id = 2077 then
	sram_write <= x"07DC0038";
end if;
if first_state_sram_input_id = 2078 then
	sram_write <= x"820020A0";
end if;
if first_state_sram_input_id = 2079 then
	sram_write <= x"02400001";
end if;
if first_state_sram_input_id = 2080 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2081 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 2082 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 2083 then
	sram_write <= x"03DC0038";
end if;
if first_state_sram_input_id = 2084 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2085 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2086 then
	sram_write <= x"8200084C";
end if;
if first_state_sram_input_id = 2087 then
	sram_write <= x"07DC0038";
end if;
if first_state_sram_input_id = 2088 then
	sram_write <= x"820020C8";
end if;
if first_state_sram_input_id = 2089 then
	sram_write <= x"0240FFFF";
end if;
if first_state_sram_input_id = 2090 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2091 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 2092 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 2093 then
	sram_write <= x"03DC0038";
end if;
if first_state_sram_input_id = 2094 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2095 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2096 then
	sram_write <= x"8200084C";
end if;
if first_state_sram_input_id = 2097 then
	sram_write <= x"07DC0038";
end if;
if first_state_sram_input_id = 2098 then
	sram_write <= x"C03C0010";
end if;
if first_state_sram_input_id = 2099 then
	sram_write <= x"C8420008";
end if;
if first_state_sram_input_id = 2100 then
	sram_write <= x"C87C0008";
end if;
if first_state_sram_input_id = 2101 then
	sram_write <= x"CC3C0030";
end if;
if first_state_sram_input_id = 2102 then
	sram_write <= x"8E462100";
end if;
if first_state_sram_input_id = 2103 then
	sram_write <= x"44446000";
end if;
if first_state_sram_input_id = 2104 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2105 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 2106 then
	sram_write <= x"03DC0040";
end if;
if first_state_sram_input_id = 2107 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2108 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2109 then
	sram_write <= x"82001270";
end if;
if first_state_sram_input_id = 2110 then
	sram_write <= x"07DC0040";
end if;
if first_state_sram_input_id = 2111 then
	sram_write <= x"8200217C";
end if;
if first_state_sram_input_id = 2112 then
	sram_write <= x"8E042158";
end if;
if first_state_sram_input_id = 2113 then
	sram_write <= x"C8800090";
end if;
if first_state_sram_input_id = 2114 then
	sram_write <= x"8E842130";
end if;
if first_state_sram_input_id = 2115 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 2116 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2117 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 2118 then
	sram_write <= x"03DC0040";
end if;
if first_state_sram_input_id = 2119 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2120 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2121 then
	sram_write <= x"82001270";
end if;
if first_state_sram_input_id = 2122 then
	sram_write <= x"07DC0040";
end if;
if first_state_sram_input_id = 2123 then
	sram_write <= x"82002154";
end if;
if first_state_sram_input_id = 2124 then
	sram_write <= x"02400001";
end if;
if first_state_sram_input_id = 2125 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2126 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 2127 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 2128 then
	sram_write <= x"03DC0040";
end if;
if first_state_sram_input_id = 2129 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2130 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2131 then
	sram_write <= x"82000B88";
end if;
if first_state_sram_input_id = 2132 then
	sram_write <= x"07DC0040";
end if;
if first_state_sram_input_id = 2133 then
	sram_write <= x"8200217C";
end if;
if first_state_sram_input_id = 2134 then
	sram_write <= x"0240FFFF";
end if;
if first_state_sram_input_id = 2135 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2136 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 2137 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 2138 then
	sram_write <= x"03DC0040";
end if;
if first_state_sram_input_id = 2139 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2140 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2141 then
	sram_write <= x"82000B88";
end if;
if first_state_sram_input_id = 2142 then
	sram_write <= x"07DC0040";
end if;
if first_state_sram_input_id = 2143 then
	sram_write <= x"C03C0010";
end if;
if first_state_sram_input_id = 2144 then
	sram_write <= x"C8420008";
end if;
if first_state_sram_input_id = 2145 then
	sram_write <= x"C87C0008";
end if;
if first_state_sram_input_id = 2146 then
	sram_write <= x"CC3C0038";
end if;
if first_state_sram_input_id = 2147 then
	sram_write <= x"8E4621B4";
end if;
if first_state_sram_input_id = 2148 then
	sram_write <= x"44446000";
end if;
if first_state_sram_input_id = 2149 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2150 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 2151 then
	sram_write <= x"03DC0048";
end if;
if first_state_sram_input_id = 2152 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2153 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2154 then
	sram_write <= x"82000EC4";
end if;
if first_state_sram_input_id = 2155 then
	sram_write <= x"07DC0048";
end if;
if first_state_sram_input_id = 2156 then
	sram_write <= x"82002230";
end if;
if first_state_sram_input_id = 2157 then
	sram_write <= x"8E04220C";
end if;
if first_state_sram_input_id = 2158 then
	sram_write <= x"C8800090";
end if;
if first_state_sram_input_id = 2159 then
	sram_write <= x"8E8421E4";
end if;
if first_state_sram_input_id = 2160 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 2161 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2162 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 2163 then
	sram_write <= x"03DC0048";
end if;
if first_state_sram_input_id = 2164 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2165 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2166 then
	sram_write <= x"82000EC4";
end if;
if first_state_sram_input_id = 2167 then
	sram_write <= x"07DC0048";
end if;
if first_state_sram_input_id = 2168 then
	sram_write <= x"82002208";
end if;
if first_state_sram_input_id = 2169 then
	sram_write <= x"02400001";
end if;
if first_state_sram_input_id = 2170 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2171 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 2172 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 2173 then
	sram_write <= x"03DC0048";
end if;
if first_state_sram_input_id = 2174 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2175 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2176 then
	sram_write <= x"8200084C";
end if;
if first_state_sram_input_id = 2177 then
	sram_write <= x"07DC0048";
end if;
if first_state_sram_input_id = 2178 then
	sram_write <= x"82002230";
end if;
if first_state_sram_input_id = 2179 then
	sram_write <= x"0240FFFF";
end if;
if first_state_sram_input_id = 2180 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2181 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 2182 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 2183 then
	sram_write <= x"03DC0048";
end if;
if first_state_sram_input_id = 2184 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2185 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2186 then
	sram_write <= x"8200084C";
end if;
if first_state_sram_input_id = 2187 then
	sram_write <= x"07DC0048";
end if;
if first_state_sram_input_id = 2188 then
	sram_write <= x"C85C0038";
end if;
if first_state_sram_input_id = 2189 then
	sram_write <= x"C87C0028";
end if;
if first_state_sram_input_id = 2190 then
	sram_write <= x"48864000";
end if;
if first_state_sram_input_id = 2191 then
	sram_write <= x"C8BC0030";
end if;
if first_state_sram_input_id = 2192 then
	sram_write <= x"C8DC0020";
end if;
if first_state_sram_input_id = 2193 then
	sram_write <= x"48ECA000";
end if;
if first_state_sram_input_id = 2194 then
	sram_write <= x"490E4000";
end if;
if first_state_sram_input_id = 2195 then
	sram_write <= x"C93C0018";
end if;
if first_state_sram_input_id = 2196 then
	sram_write <= x"49522000";
end if;
if first_state_sram_input_id = 2197 then
	sram_write <= x"45114000";
end if;
if first_state_sram_input_id = 2198 then
	sram_write <= x"4952A000";
end if;
if first_state_sram_input_id = 2199 then
	sram_write <= x"49744000";
end if;
if first_state_sram_input_id = 2200 then
	sram_write <= x"498C2000";
end if;
if first_state_sram_input_id = 2201 then
	sram_write <= x"41778000";
end if;
if first_state_sram_input_id = 2202 then
	sram_write <= x"49862000";
end if;
if first_state_sram_input_id = 2203 then
	sram_write <= x"48EE2000";
end if;
if first_state_sram_input_id = 2204 then
	sram_write <= x"49B24000";
end if;
if first_state_sram_input_id = 2205 then
	sram_write <= x"40EFA000";
end if;
if first_state_sram_input_id = 2206 then
	sram_write <= x"48342000";
end if;
if first_state_sram_input_id = 2207 then
	sram_write <= x"484C4000";
end if;
if first_state_sram_input_id = 2208 then
	sram_write <= x"44224000";
end if;
if first_state_sram_input_id = 2209 then
	sram_write <= x"4440A000";
end if;
if first_state_sram_input_id = 2210 then
	sram_write <= x"48AC6000";
end if;
if first_state_sram_input_id = 2211 then
	sram_write <= x"48726000";
end if;
if first_state_sram_input_id = 2212 then
	sram_write <= x"C03C0000";
end if;
if first_state_sram_input_id = 2213 then
	sram_write <= x"C8C20000";
end if;
if first_state_sram_input_id = 2214 then
	sram_write <= x"C9220004";
end if;
if first_state_sram_input_id = 2215 then
	sram_write <= x"C9420008";
end if;
if first_state_sram_input_id = 2216 then
	sram_write <= x"49A88000";
end if;
if first_state_sram_input_id = 2217 then
	sram_write <= x"49ADA000";
end if;
if first_state_sram_input_id = 2218 then
	sram_write <= x"49D98000";
end if;
if first_state_sram_input_id = 2219 then
	sram_write <= x"49D3C000";
end if;
if first_state_sram_input_id = 2220 then
	sram_write <= x"41BBC000";
end if;
if first_state_sram_input_id = 2221 then
	sram_write <= x"49C44000";
end if;
if first_state_sram_input_id = 2222 then
	sram_write <= x"49D5C000";
end if;
if first_state_sram_input_id = 2223 then
	sram_write <= x"41BBC000";
end if;
if first_state_sram_input_id = 2224 then
	sram_write <= x"CDA20000";
end if;
if first_state_sram_input_id = 2225 then
	sram_write <= x"49B10000";
end if;
if first_state_sram_input_id = 2226 then
	sram_write <= x"49ADA000";
end if;
if first_state_sram_input_id = 2227 then
	sram_write <= x"49CEE000";
end if;
if first_state_sram_input_id = 2228 then
	sram_write <= x"49D3C000";
end if;
if first_state_sram_input_id = 2229 then
	sram_write <= x"41BBC000";
end if;
if first_state_sram_input_id = 2230 then
	sram_write <= x"49CAA000";
end if;
if first_state_sram_input_id = 2231 then
	sram_write <= x"49D5C000";
end if;
if first_state_sram_input_id = 2232 then
	sram_write <= x"41BBC000";
end if;
if first_state_sram_input_id = 2233 then
	sram_write <= x"CDA20004";
end if;
if first_state_sram_input_id = 2234 then
	sram_write <= x"49B76000";
end if;
if first_state_sram_input_id = 2235 then
	sram_write <= x"49ADA000";
end if;
if first_state_sram_input_id = 2236 then
	sram_write <= x"49C22000";
end if;
if first_state_sram_input_id = 2237 then
	sram_write <= x"49D3C000";
end if;
if first_state_sram_input_id = 2238 then
	sram_write <= x"41BBC000";
end if;
if first_state_sram_input_id = 2239 then
	sram_write <= x"49C66000";
end if;
if first_state_sram_input_id = 2240 then
	sram_write <= x"49D5C000";
end if;
if first_state_sram_input_id = 2241 then
	sram_write <= x"41BBC000";
end if;
if first_state_sram_input_id = 2242 then
	sram_write <= x"CDA20008";
end if;
if first_state_sram_input_id = 2243 then
	sram_write <= x"C9A00080";
end if;
if first_state_sram_input_id = 2244 then
	sram_write <= x"49CD0000";
end if;
if first_state_sram_input_id = 2245 then
	sram_write <= x"49DD6000";
end if;
if first_state_sram_input_id = 2246 then
	sram_write <= x"49F2E000";
end if;
if first_state_sram_input_id = 2247 then
	sram_write <= x"49FE2000";
end if;
if first_state_sram_input_id = 2248 then
	sram_write <= x"41DDE000";
end if;
if first_state_sram_input_id = 2249 then
	sram_write <= x"49F4A000";
end if;
if first_state_sram_input_id = 2250 then
	sram_write <= x"49FE6000";
end if;
if first_state_sram_input_id = 2251 then
	sram_write <= x"41DDE000";
end if;
if first_state_sram_input_id = 2252 then
	sram_write <= x"49DBC000";
end if;
if first_state_sram_input_id = 2253 then
	sram_write <= x"C03C0010";
end if;
if first_state_sram_input_id = 2254 then
	sram_write <= x"CDC20000";
end if;
if first_state_sram_input_id = 2255 then
	sram_write <= x"488C8000";
end if;
if first_state_sram_input_id = 2256 then
	sram_write <= x"48C96000";
end if;
if first_state_sram_input_id = 2257 then
	sram_write <= x"49338000";
end if;
if first_state_sram_input_id = 2258 then
	sram_write <= x"48322000";
end if;
if first_state_sram_input_id = 2259 then
	sram_write <= x"402C2000";
end if;
if first_state_sram_input_id = 2260 then
	sram_write <= x"48544000";
end if;
if first_state_sram_input_id = 2261 then
	sram_write <= x"48646000";
end if;
if first_state_sram_input_id = 2262 then
	sram_write <= x"40226000";
end if;
if first_state_sram_input_id = 2263 then
	sram_write <= x"483A2000";
end if;
if first_state_sram_input_id = 2264 then
	sram_write <= x"CC220004";
end if;
if first_state_sram_input_id = 2265 then
	sram_write <= x"48290000";
end if;
if first_state_sram_input_id = 2266 then
	sram_write <= x"4872E000";
end if;
if first_state_sram_input_id = 2267 then
	sram_write <= x"40226000";
end if;
if first_state_sram_input_id = 2268 then
	sram_write <= x"4844A000";
end if;
if first_state_sram_input_id = 2269 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 2270 then
	sram_write <= x"483A2000";
end if;
if first_state_sram_input_id = 2271 then
	sram_write <= x"CC220008";
end if;
if first_state_sram_input_id = 2272 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 2273 then
	sram_write <= x"C43C0000";
end if;
if first_state_sram_input_id = 2274 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2275 then
	sram_write <= x"03DC000C";
end if;
if first_state_sram_input_id = 2276 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2277 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2278 then
	sram_write <= x"82000794";
end if;
if first_state_sram_input_id = 2279 then
	sram_write <= x"07DC000C";
end if;
if first_state_sram_input_id = 2280 then
	sram_write <= x"0240FFFF";
end if;
if first_state_sram_input_id = 2281 then
	sram_write <= x"82242928";
end if;
if first_state_sram_input_id = 2282 then
	sram_write <= x"C43C0004";
end if;
if first_state_sram_input_id = 2283 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2284 then
	sram_write <= x"03DC0010";
end if;
if first_state_sram_input_id = 2285 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2286 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2287 then
	sram_write <= x"82000794";
end if;
if first_state_sram_input_id = 2288 then
	sram_write <= x"07DC0010";
end if;
if first_state_sram_input_id = 2289 then
	sram_write <= x"C43C0008";
end if;
if first_state_sram_input_id = 2290 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2291 then
	sram_write <= x"03DC0014";
end if;
if first_state_sram_input_id = 2292 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2293 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2294 then
	sram_write <= x"82000794";
end if;
if first_state_sram_input_id = 2295 then
	sram_write <= x"07DC0014";
end if;
if first_state_sram_input_id = 2296 then
	sram_write <= x"C43C000C";
end if;
if first_state_sram_input_id = 2297 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2298 then
	sram_write <= x"03DC0018";
end if;
if first_state_sram_input_id = 2299 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2300 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2301 then
	sram_write <= x"82000794";
end if;
if first_state_sram_input_id = 2302 then
	sram_write <= x"07DC0018";
end if;
if first_state_sram_input_id = 2303 then
	sram_write <= x"02400003";
end if;
if first_state_sram_input_id = 2304 then
	sram_write <= x"40200000";
end if;
if first_state_sram_input_id = 2305 then
	sram_write <= x"C43C0010";
end if;
if first_state_sram_input_id = 2306 then
	sram_write <= x"CC3C0018";
end if;
if first_state_sram_input_id = 2307 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2308 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 2309 then
	sram_write <= x"03DC0028";
end if;
if first_state_sram_input_id = 2310 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2311 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2312 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 2313 then
	sram_write <= x"07DC0028";
end if;
if first_state_sram_input_id = 2314 then
	sram_write <= x"C43C0020";
end if;
if first_state_sram_input_id = 2315 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2316 then
	sram_write <= x"03DC002C";
end if;
if first_state_sram_input_id = 2317 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2318 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2319 then
	sram_write <= x"820007C0";
end if;
if first_state_sram_input_id = 2320 then
	sram_write <= x"07DC002C";
end if;
if first_state_sram_input_id = 2321 then
	sram_write <= x"C03C0020";
end if;
if first_state_sram_input_id = 2322 then
	sram_write <= x"CC220000";
end if;
if first_state_sram_input_id = 2323 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2324 then
	sram_write <= x"03DC002C";
end if;
if first_state_sram_input_id = 2325 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2326 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2327 then
	sram_write <= x"820007C0";
end if;
if first_state_sram_input_id = 2328 then
	sram_write <= x"07DC002C";
end if;
if first_state_sram_input_id = 2329 then
	sram_write <= x"C03C0020";
end if;
if first_state_sram_input_id = 2330 then
	sram_write <= x"CC220004";
end if;
if first_state_sram_input_id = 2331 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2332 then
	sram_write <= x"03DC002C";
end if;
if first_state_sram_input_id = 2333 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2334 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2335 then
	sram_write <= x"820007C0";
end if;
if first_state_sram_input_id = 2336 then
	sram_write <= x"07DC002C";
end if;
if first_state_sram_input_id = 2337 then
	sram_write <= x"C03C0020";
end if;
if first_state_sram_input_id = 2338 then
	sram_write <= x"CC220008";
end if;
if first_state_sram_input_id = 2339 then
	sram_write <= x"02400003";
end if;
if first_state_sram_input_id = 2340 then
	sram_write <= x"C83C0018";
end if;
if first_state_sram_input_id = 2341 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2342 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 2343 then
	sram_write <= x"03DC002C";
end if;
if first_state_sram_input_id = 2344 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2345 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2346 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 2347 then
	sram_write <= x"07DC002C";
end if;
if first_state_sram_input_id = 2348 then
	sram_write <= x"C43C0024";
end if;
if first_state_sram_input_id = 2349 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2350 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 2351 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2352 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2353 then
	sram_write <= x"820007C0";
end if;
if first_state_sram_input_id = 2354 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 2355 then
	sram_write <= x"C03C0024";
end if;
if first_state_sram_input_id = 2356 then
	sram_write <= x"CC220000";
end if;
if first_state_sram_input_id = 2357 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2358 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 2359 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2360 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2361 then
	sram_write <= x"820007C0";
end if;
if first_state_sram_input_id = 2362 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 2363 then
	sram_write <= x"C03C0024";
end if;
if first_state_sram_input_id = 2364 then
	sram_write <= x"CC220004";
end if;
if first_state_sram_input_id = 2365 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2366 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 2367 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2368 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2369 then
	sram_write <= x"820007C0";
end if;
if first_state_sram_input_id = 2370 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 2371 then
	sram_write <= x"C03C0024";
end if;
if first_state_sram_input_id = 2372 then
	sram_write <= x"CC220008";
end if;
if first_state_sram_input_id = 2373 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2374 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 2375 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2376 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2377 then
	sram_write <= x"820007C0";
end if;
if first_state_sram_input_id = 2378 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 2379 then
	sram_write <= x"8E202538";
end if;
if first_state_sram_input_id = 2380 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 2381 then
	sram_write <= x"8200253C";
end if;
if first_state_sram_input_id = 2382 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 2383 then
	sram_write <= x"02400002";
end if;
if first_state_sram_input_id = 2384 then
	sram_write <= x"C85C0018";
end if;
if first_state_sram_input_id = 2385 then
	sram_write <= x"CC3C0028";
end if;
if first_state_sram_input_id = 2386 then
	sram_write <= x"C43C0030";
end if;
if first_state_sram_input_id = 2387 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2388 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 2389 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 2390 then
	sram_write <= x"03DC003C";
end if;
if first_state_sram_input_id = 2391 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2392 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2393 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 2394 then
	sram_write <= x"07DC003C";
end if;
if first_state_sram_input_id = 2395 then
	sram_write <= x"C43C0034";
end if;
if first_state_sram_input_id = 2396 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2397 then
	sram_write <= x"03DC0040";
end if;
if first_state_sram_input_id = 2398 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2399 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2400 then
	sram_write <= x"820007C0";
end if;
if first_state_sram_input_id = 2401 then
	sram_write <= x"07DC0040";
end if;
if first_state_sram_input_id = 2402 then
	sram_write <= x"C03C0034";
end if;
if first_state_sram_input_id = 2403 then
	sram_write <= x"CC220000";
end if;
if first_state_sram_input_id = 2404 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2405 then
	sram_write <= x"03DC0040";
end if;
if first_state_sram_input_id = 2406 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2407 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2408 then
	sram_write <= x"820007C0";
end if;
if first_state_sram_input_id = 2409 then
	sram_write <= x"07DC0040";
end if;
if first_state_sram_input_id = 2410 then
	sram_write <= x"C03C0034";
end if;
if first_state_sram_input_id = 2411 then
	sram_write <= x"CC220004";
end if;
if first_state_sram_input_id = 2412 then
	sram_write <= x"02400003";
end if;
if first_state_sram_input_id = 2413 then
	sram_write <= x"C83C0018";
end if;
if first_state_sram_input_id = 2414 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2415 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 2416 then
	sram_write <= x"03DC0040";
end if;
if first_state_sram_input_id = 2417 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2418 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2419 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 2420 then
	sram_write <= x"07DC0040";
end if;
if first_state_sram_input_id = 2421 then
	sram_write <= x"C43C0038";
end if;
if first_state_sram_input_id = 2422 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2423 then
	sram_write <= x"03DC0044";
end if;
if first_state_sram_input_id = 2424 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2425 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2426 then
	sram_write <= x"820007C0";
end if;
if first_state_sram_input_id = 2427 then
	sram_write <= x"07DC0044";
end if;
if first_state_sram_input_id = 2428 then
	sram_write <= x"C03C0038";
end if;
if first_state_sram_input_id = 2429 then
	sram_write <= x"CC220000";
end if;
if first_state_sram_input_id = 2430 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2431 then
	sram_write <= x"03DC0044";
end if;
if first_state_sram_input_id = 2432 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2433 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2434 then
	sram_write <= x"820007C0";
end if;
if first_state_sram_input_id = 2435 then
	sram_write <= x"07DC0044";
end if;
if first_state_sram_input_id = 2436 then
	sram_write <= x"C03C0038";
end if;
if first_state_sram_input_id = 2437 then
	sram_write <= x"CC220004";
end if;
if first_state_sram_input_id = 2438 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2439 then
	sram_write <= x"03DC0044";
end if;
if first_state_sram_input_id = 2440 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2441 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2442 then
	sram_write <= x"820007C0";
end if;
if first_state_sram_input_id = 2443 then
	sram_write <= x"07DC0044";
end if;
if first_state_sram_input_id = 2444 then
	sram_write <= x"C03C0038";
end if;
if first_state_sram_input_id = 2445 then
	sram_write <= x"CC220008";
end if;
if first_state_sram_input_id = 2446 then
	sram_write <= x"02400003";
end if;
if first_state_sram_input_id = 2447 then
	sram_write <= x"C83C0018";
end if;
if first_state_sram_input_id = 2448 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2449 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 2450 then
	sram_write <= x"03DC0044";
end if;
if first_state_sram_input_id = 2451 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2452 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2453 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 2454 then
	sram_write <= x"07DC0044";
end if;
if first_state_sram_input_id = 2455 then
	sram_write <= x"C05C0010";
end if;
if first_state_sram_input_id = 2456 then
	sram_write <= x"824026E8";
end if;
if first_state_sram_input_id = 2457 then
	sram_write <= x"C43C003C";
end if;
if first_state_sram_input_id = 2458 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2459 then
	sram_write <= x"03DC0048";
end if;
if first_state_sram_input_id = 2460 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2461 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2462 then
	sram_write <= x"820007C0";
end if;
if first_state_sram_input_id = 2463 then
	sram_write <= x"07DC0048";
end if;
if first_state_sram_input_id = 2464 then
	sram_write <= x"C840008C";
end if;
if first_state_sram_input_id = 2465 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 2466 then
	sram_write <= x"C03C003C";
end if;
if first_state_sram_input_id = 2467 then
	sram_write <= x"CC220000";
end if;
if first_state_sram_input_id = 2468 then
	sram_write <= x"CC5C0040";
end if;
if first_state_sram_input_id = 2469 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2470 then
	sram_write <= x"03DC0050";
end if;
if first_state_sram_input_id = 2471 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2472 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2473 then
	sram_write <= x"820007C0";
end if;
if first_state_sram_input_id = 2474 then
	sram_write <= x"07DC0050";
end if;
if first_state_sram_input_id = 2475 then
	sram_write <= x"C85C0040";
end if;
if first_state_sram_input_id = 2476 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 2477 then
	sram_write <= x"C03C003C";
end if;
if first_state_sram_input_id = 2478 then
	sram_write <= x"CC220004";
end if;
if first_state_sram_input_id = 2479 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2480 then
	sram_write <= x"03DC0050";
end if;
if first_state_sram_input_id = 2481 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2482 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2483 then
	sram_write <= x"820007C0";
end if;
if first_state_sram_input_id = 2484 then
	sram_write <= x"07DC0050";
end if;
if first_state_sram_input_id = 2485 then
	sram_write <= x"C85C0040";
end if;
if first_state_sram_input_id = 2486 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 2487 then
	sram_write <= x"C03C003C";
end if;
if first_state_sram_input_id = 2488 then
	sram_write <= x"CC220008";
end if;
if first_state_sram_input_id = 2489 then
	sram_write <= x"820026E8";
end if;
if first_state_sram_input_id = 2490 then
	sram_write <= x"02400002";
end if;
if first_state_sram_input_id = 2491 then
	sram_write <= x"C07C0008";
end if;
if first_state_sram_input_id = 2492 then
	sram_write <= x"826426FC";
end if;
if first_state_sram_input_id = 2493 then
	sram_write <= x"C05C0030";
end if;
if first_state_sram_input_id = 2494 then
	sram_write <= x"82002700";
end if;
if first_state_sram_input_id = 2495 then
	sram_write <= x"02400001";
end if;
if first_state_sram_input_id = 2496 then
	sram_write <= x"02800004";
end if;
if first_state_sram_input_id = 2497 then
	sram_write <= x"C83C0018";
end if;
if first_state_sram_input_id = 2498 then
	sram_write <= x"C45C0048";
end if;
if first_state_sram_input_id = 2499 then
	sram_write <= x"C43C003C";
end if;
if first_state_sram_input_id = 2500 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2501 then
	sram_write <= x"00280000";
end if;
if first_state_sram_input_id = 2502 then
	sram_write <= x"03DC0054";
end if;
if first_state_sram_input_id = 2503 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2504 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2505 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 2506 then
	sram_write <= x"07DC0054";
end if;
if first_state_sram_input_id = 2507 then
	sram_write <= x"005A0000";
end if;
if first_state_sram_input_id = 2508 then
	sram_write <= x"03BA002C";
end if;
if first_state_sram_input_id = 2509 then
	sram_write <= x"C4240028";
end if;
if first_state_sram_input_id = 2510 then
	sram_write <= x"C03C003C";
end if;
if first_state_sram_input_id = 2511 then
	sram_write <= x"C4240024";
end if;
if first_state_sram_input_id = 2512 then
	sram_write <= x"C07C0038";
end if;
if first_state_sram_input_id = 2513 then
	sram_write <= x"C4640020";
end if;
if first_state_sram_input_id = 2514 then
	sram_write <= x"C07C0034";
end if;
if first_state_sram_input_id = 2515 then
	sram_write <= x"C464001C";
end if;
if first_state_sram_input_id = 2516 then
	sram_write <= x"C07C0048";
end if;
if first_state_sram_input_id = 2517 then
	sram_write <= x"C4640018";
end if;
if first_state_sram_input_id = 2518 then
	sram_write <= x"C07C0024";
end if;
if first_state_sram_input_id = 2519 then
	sram_write <= x"C4640014";
end if;
if first_state_sram_input_id = 2520 then
	sram_write <= x"C07C0020";
end if;
if first_state_sram_input_id = 2521 then
	sram_write <= x"C4640010";
end if;
if first_state_sram_input_id = 2522 then
	sram_write <= x"C09C0010";
end if;
if first_state_sram_input_id = 2523 then
	sram_write <= x"C484000C";
end if;
if first_state_sram_input_id = 2524 then
	sram_write <= x"C0BC000C";
end if;
if first_state_sram_input_id = 2525 then
	sram_write <= x"C4A40008";
end if;
if first_state_sram_input_id = 2526 then
	sram_write <= x"C0BC0008";
end if;
if first_state_sram_input_id = 2527 then
	sram_write <= x"C4A40004";
end if;
if first_state_sram_input_id = 2528 then
	sram_write <= x"C0DC0004";
end if;
if first_state_sram_input_id = 2529 then
	sram_write <= x"C4C40000";
end if;
if first_state_sram_input_id = 2530 then
	sram_write <= x"02C000C8";
end if;
if first_state_sram_input_id = 2531 then
	sram_write <= x"C0FC0000";
end if;
if first_state_sram_input_id = 2532 then
	sram_write <= x"22EE0220";
end if;
if first_state_sram_input_id = 2533 then
	sram_write <= x"D44CE000";
end if;
if first_state_sram_input_id = 2534 then
	sram_write <= x"02400003";
end if;
if first_state_sram_input_id = 2535 then
	sram_write <= x"82A427E0";
end if;
if first_state_sram_input_id = 2536 then
	sram_write <= x"02400002";
end if;
if first_state_sram_input_id = 2537 then
	sram_write <= x"82A427AC";
end if;
if first_state_sram_input_id = 2538 then
	sram_write <= x"820027DC";
end if;
if first_state_sram_input_id = 2539 then
	sram_write <= x"C83C0028";
end if;
if first_state_sram_input_id = 2540 then
	sram_write <= x"8E2027BC";
end if;
if first_state_sram_input_id = 2541 then
	sram_write <= x"02400001";
end if;
if first_state_sram_input_id = 2542 then
	sram_write <= x"820027C0";
end if;
if first_state_sram_input_id = 2543 then
	sram_write <= x"02400000";
end if;
if first_state_sram_input_id = 2544 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2545 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 2546 then
	sram_write <= x"03DC0054";
end if;
if first_state_sram_input_id = 2547 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2548 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2549 then
	sram_write <= x"8200161C";
end if;
if first_state_sram_input_id = 2550 then
	sram_write <= x"07DC0054";
end if;
if first_state_sram_input_id = 2551 then
	sram_write <= x"820028F4";
end if;
if first_state_sram_input_id = 2552 then
	sram_write <= x"C8260000";
end if;
if first_state_sram_input_id = 2553 then
	sram_write <= x"8A202830";
end if;
if first_state_sram_input_id = 2554 then
	sram_write <= x"8A202800";
end if;
if first_state_sram_input_id = 2555 then
	sram_write <= x"8E0227F8";
end if;
if first_state_sram_input_id = 2556 then
	sram_write <= x"C840007C";
end if;
if first_state_sram_input_id = 2557 then
	sram_write <= x"820027FC";
end if;
if first_state_sram_input_id = 2558 then
	sram_write <= x"C84000A8";
end if;
if first_state_sram_input_id = 2559 then
	sram_write <= x"82002804";
end if;
if first_state_sram_input_id = 2560 then
	sram_write <= x"40400000";
end if;
if first_state_sram_input_id = 2561 then
	sram_write <= x"48222000";
end if;
if first_state_sram_input_id = 2562 then
	sram_write <= x"CC5C0050";
end if;
if first_state_sram_input_id = 2563 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2564 then
	sram_write <= x"03DC0060";
end if;
if first_state_sram_input_id = 2565 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2566 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2567 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 2568 then
	sram_write <= x"07DC0060";
end if;
if first_state_sram_input_id = 2569 then
	sram_write <= x"C85C0050";
end if;
if first_state_sram_input_id = 2570 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 2571 then
	sram_write <= x"82002834";
end if;
if first_state_sram_input_id = 2572 then
	sram_write <= x"40200000";
end if;
if first_state_sram_input_id = 2573 then
	sram_write <= x"C03C0020";
end if;
if first_state_sram_input_id = 2574 then
	sram_write <= x"CC220000";
end if;
if first_state_sram_input_id = 2575 then
	sram_write <= x"C8220004";
end if;
if first_state_sram_input_id = 2576 then
	sram_write <= x"8A20288C";
end if;
if first_state_sram_input_id = 2577 then
	sram_write <= x"8A20285C";
end if;
if first_state_sram_input_id = 2578 then
	sram_write <= x"8E022854";
end if;
if first_state_sram_input_id = 2579 then
	sram_write <= x"C840007C";
end if;
if first_state_sram_input_id = 2580 then
	sram_write <= x"82002858";
end if;
if first_state_sram_input_id = 2581 then
	sram_write <= x"C84000A8";
end if;
if first_state_sram_input_id = 2582 then
	sram_write <= x"82002860";
end if;
if first_state_sram_input_id = 2583 then
	sram_write <= x"40400000";
end if;
if first_state_sram_input_id = 2584 then
	sram_write <= x"48222000";
end if;
if first_state_sram_input_id = 2585 then
	sram_write <= x"CC5C0058";
end if;
if first_state_sram_input_id = 2586 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2587 then
	sram_write <= x"03DC0068";
end if;
if first_state_sram_input_id = 2588 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2589 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2590 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 2591 then
	sram_write <= x"07DC0068";
end if;
if first_state_sram_input_id = 2592 then
	sram_write <= x"C85C0058";
end if;
if first_state_sram_input_id = 2593 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 2594 then
	sram_write <= x"82002890";
end if;
if first_state_sram_input_id = 2595 then
	sram_write <= x"40200000";
end if;
if first_state_sram_input_id = 2596 then
	sram_write <= x"C03C0020";
end if;
if first_state_sram_input_id = 2597 then
	sram_write <= x"CC220004";
end if;
if first_state_sram_input_id = 2598 then
	sram_write <= x"C8220008";
end if;
if first_state_sram_input_id = 2599 then
	sram_write <= x"8A2028E8";
end if;
if first_state_sram_input_id = 2600 then
	sram_write <= x"8A2028B8";
end if;
if first_state_sram_input_id = 2601 then
	sram_write <= x"8E0228B0";
end if;
if first_state_sram_input_id = 2602 then
	sram_write <= x"C840007C";
end if;
if first_state_sram_input_id = 2603 then
	sram_write <= x"820028B4";
end if;
if first_state_sram_input_id = 2604 then
	sram_write <= x"C84000A8";
end if;
if first_state_sram_input_id = 2605 then
	sram_write <= x"820028BC";
end if;
if first_state_sram_input_id = 2606 then
	sram_write <= x"40400000";
end if;
if first_state_sram_input_id = 2607 then
	sram_write <= x"48222000";
end if;
if first_state_sram_input_id = 2608 then
	sram_write <= x"CC5C0060";
end if;
if first_state_sram_input_id = 2609 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2610 then
	sram_write <= x"03DC0070";
end if;
if first_state_sram_input_id = 2611 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2612 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2613 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 2614 then
	sram_write <= x"07DC0070";
end if;
if first_state_sram_input_id = 2615 then
	sram_write <= x"C85C0060";
end if;
if first_state_sram_input_id = 2616 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 2617 then
	sram_write <= x"820028EC";
end if;
if first_state_sram_input_id = 2618 then
	sram_write <= x"40200000";
end if;
if first_state_sram_input_id = 2619 then
	sram_write <= x"C03C0020";
end if;
if first_state_sram_input_id = 2620 then
	sram_write <= x"CC220008";
end if;
if first_state_sram_input_id = 2621 then
	sram_write <= x"C03C0010";
end if;
if first_state_sram_input_id = 2622 then
	sram_write <= x"82202920";
end if;
if first_state_sram_input_id = 2623 then
	sram_write <= x"C03C0020";
end if;
if first_state_sram_input_id = 2624 then
	sram_write <= x"C05C003C";
end if;
if first_state_sram_input_id = 2625 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2626 then
	sram_write <= x"03DC0070";
end if;
if first_state_sram_input_id = 2627 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2628 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2629 then
	sram_write <= x"82001E04";
end if;
if first_state_sram_input_id = 2630 then
	sram_write <= x"07DC0070";
end if;
if first_state_sram_input_id = 2631 then
	sram_write <= x"82002920";
end if;
if first_state_sram_input_id = 2632 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 2633 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 2634 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 2635 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 2636 then
	sram_write <= x"0240003C";
end if;
if first_state_sram_input_id = 2637 then
	sram_write <= x"8624293C";
end if;
if first_state_sram_input_id = 2638 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 2639 then
	sram_write <= x"C43C0000";
end if;
if first_state_sram_input_id = 2640 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2641 then
	sram_write <= x"03DC000C";
end if;
if first_state_sram_input_id = 2642 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2643 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2644 then
	sram_write <= x"82002384";
end if;
if first_state_sram_input_id = 2645 then
	sram_write <= x"07DC000C";
end if;
if first_state_sram_input_id = 2646 then
	sram_write <= x"82202A34";
end if;
if first_state_sram_input_id = 2647 then
	sram_write <= x"C03C0000";
end if;
if first_state_sram_input_id = 2648 then
	sram_write <= x"02220001";
end if;
if first_state_sram_input_id = 2649 then
	sram_write <= x"0240003C";
end if;
if first_state_sram_input_id = 2650 then
	sram_write <= x"86242970";
end if;
if first_state_sram_input_id = 2651 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 2652 then
	sram_write <= x"C43C0004";
end if;
if first_state_sram_input_id = 2653 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2654 then
	sram_write <= x"03DC0010";
end if;
if first_state_sram_input_id = 2655 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2656 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2657 then
	sram_write <= x"82002384";
end if;
if first_state_sram_input_id = 2658 then
	sram_write <= x"07DC0010";
end if;
if first_state_sram_input_id = 2659 then
	sram_write <= x"82202A24";
end if;
if first_state_sram_input_id = 2660 then
	sram_write <= x"C03C0004";
end if;
if first_state_sram_input_id = 2661 then
	sram_write <= x"02220001";
end if;
if first_state_sram_input_id = 2662 then
	sram_write <= x"0240003C";
end if;
if first_state_sram_input_id = 2663 then
	sram_write <= x"862429A4";
end if;
if first_state_sram_input_id = 2664 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 2665 then
	sram_write <= x"C43C0008";
end if;
if first_state_sram_input_id = 2666 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2667 then
	sram_write <= x"03DC0014";
end if;
if first_state_sram_input_id = 2668 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2669 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2670 then
	sram_write <= x"82002384";
end if;
if first_state_sram_input_id = 2671 then
	sram_write <= x"07DC0014";
end if;
if first_state_sram_input_id = 2672 then
	sram_write <= x"82202A14";
end if;
if first_state_sram_input_id = 2673 then
	sram_write <= x"C03C0008";
end if;
if first_state_sram_input_id = 2674 then
	sram_write <= x"02220001";
end if;
if first_state_sram_input_id = 2675 then
	sram_write <= x"0240003C";
end if;
if first_state_sram_input_id = 2676 then
	sram_write <= x"862429D8";
end if;
if first_state_sram_input_id = 2677 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 2678 then
	sram_write <= x"C43C000C";
end if;
if first_state_sram_input_id = 2679 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2680 then
	sram_write <= x"03DC0018";
end if;
if first_state_sram_input_id = 2681 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2682 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2683 then
	sram_write <= x"82002384";
end if;
if first_state_sram_input_id = 2684 then
	sram_write <= x"07DC0018";
end if;
if first_state_sram_input_id = 2685 then
	sram_write <= x"82202A04";
end if;
if first_state_sram_input_id = 2686 then
	sram_write <= x"C03C000C";
end if;
if first_state_sram_input_id = 2687 then
	sram_write <= x"02220001";
end if;
if first_state_sram_input_id = 2688 then
	sram_write <= x"82002930";
end if;
if first_state_sram_input_id = 2689 then
	sram_write <= x"022000C4";
end if;
if first_state_sram_input_id = 2690 then
	sram_write <= x"C05C000C";
end if;
if first_state_sram_input_id = 2691 then
	sram_write <= x"C4420000";
end if;
if first_state_sram_input_id = 2692 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 2693 then
	sram_write <= x"022000C4";
end if;
if first_state_sram_input_id = 2694 then
	sram_write <= x"C05C0008";
end if;
if first_state_sram_input_id = 2695 then
	sram_write <= x"C4420000";
end if;
if first_state_sram_input_id = 2696 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 2697 then
	sram_write <= x"022000C4";
end if;
if first_state_sram_input_id = 2698 then
	sram_write <= x"C05C0004";
end if;
if first_state_sram_input_id = 2699 then
	sram_write <= x"C4420000";
end if;
if first_state_sram_input_id = 2700 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 2701 then
	sram_write <= x"022000C4";
end if;
if first_state_sram_input_id = 2702 then
	sram_write <= x"C05C0000";
end if;
if first_state_sram_input_id = 2703 then
	sram_write <= x"C4420000";
end if;
if first_state_sram_input_id = 2704 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 2705 then
	sram_write <= x"C43C0000";
end if;
if first_state_sram_input_id = 2706 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2707 then
	sram_write <= x"03DC000C";
end if;
if first_state_sram_input_id = 2708 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2709 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2710 then
	sram_write <= x"82000794";
end if;
if first_state_sram_input_id = 2711 then
	sram_write <= x"07DC000C";
end if;
if first_state_sram_input_id = 2712 then
	sram_write <= x"0240FFFF";
end if;
if first_state_sram_input_id = 2713 then
	sram_write <= x"82242BDC";
end if;
if first_state_sram_input_id = 2714 then
	sram_write <= x"C05C0000";
end if;
if first_state_sram_input_id = 2715 then
	sram_write <= x"02640001";
end if;
if first_state_sram_input_id = 2716 then
	sram_write <= x"C43C0004";
end if;
if first_state_sram_input_id = 2717 then
	sram_write <= x"C47C0008";
end if;
if first_state_sram_input_id = 2718 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2719 then
	sram_write <= x"03DC0014";
end if;
if first_state_sram_input_id = 2720 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2721 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2722 then
	sram_write <= x"82000794";
end if;
if first_state_sram_input_id = 2723 then
	sram_write <= x"07DC0014";
end if;
if first_state_sram_input_id = 2724 then
	sram_write <= x"0240FFFF";
end if;
if first_state_sram_input_id = 2725 then
	sram_write <= x"82242BA4";
end if;
if first_state_sram_input_id = 2726 then
	sram_write <= x"C05C0008";
end if;
if first_state_sram_input_id = 2727 then
	sram_write <= x"02640001";
end if;
if first_state_sram_input_id = 2728 then
	sram_write <= x"C43C000C";
end if;
if first_state_sram_input_id = 2729 then
	sram_write <= x"C47C0010";
end if;
if first_state_sram_input_id = 2730 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2731 then
	sram_write <= x"03DC001C";
end if;
if first_state_sram_input_id = 2732 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2733 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2734 then
	sram_write <= x"82000794";
end if;
if first_state_sram_input_id = 2735 then
	sram_write <= x"07DC001C";
end if;
if first_state_sram_input_id = 2736 then
	sram_write <= x"0240FFFF";
end if;
if first_state_sram_input_id = 2737 then
	sram_write <= x"82242B6C";
end if;
if first_state_sram_input_id = 2738 then
	sram_write <= x"C05C0010";
end if;
if first_state_sram_input_id = 2739 then
	sram_write <= x"02640001";
end if;
if first_state_sram_input_id = 2740 then
	sram_write <= x"C43C0014";
end if;
if first_state_sram_input_id = 2741 then
	sram_write <= x"C47C0018";
end if;
if first_state_sram_input_id = 2742 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2743 then
	sram_write <= x"03DC0024";
end if;
if first_state_sram_input_id = 2744 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2745 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2746 then
	sram_write <= x"82000794";
end if;
if first_state_sram_input_id = 2747 then
	sram_write <= x"07DC0024";
end if;
if first_state_sram_input_id = 2748 then
	sram_write <= x"0240FFFF";
end if;
if first_state_sram_input_id = 2749 then
	sram_write <= x"82242B34";
end if;
if first_state_sram_input_id = 2750 then
	sram_write <= x"C05C0018";
end if;
if first_state_sram_input_id = 2751 then
	sram_write <= x"02640001";
end if;
if first_state_sram_input_id = 2752 then
	sram_write <= x"C43C001C";
end if;
if first_state_sram_input_id = 2753 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2754 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 2755 then
	sram_write <= x"03DC0028";
end if;
if first_state_sram_input_id = 2756 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2757 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2758 then
	sram_write <= x"82002A44";
end if;
if first_state_sram_input_id = 2759 then
	sram_write <= x"07DC0028";
end if;
if first_state_sram_input_id = 2760 then
	sram_write <= x"C05C0018";
end if;
if first_state_sram_input_id = 2761 then
	sram_write <= x"22440220";
end if;
if first_state_sram_input_id = 2762 then
	sram_write <= x"C07C001C";
end if;
if first_state_sram_input_id = 2763 then
	sram_write <= x"D4624000";
end if;
if first_state_sram_input_id = 2764 then
	sram_write <= x"82002B58";
end if;
if first_state_sram_input_id = 2765 then
	sram_write <= x"C03C0018";
end if;
if first_state_sram_input_id = 2766 then
	sram_write <= x"02220001";
end if;
if first_state_sram_input_id = 2767 then
	sram_write <= x"0240FFFF";
end if;
if first_state_sram_input_id = 2768 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2769 then
	sram_write <= x"03DC0028";
end if;
if first_state_sram_input_id = 2770 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2771 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2772 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 2773 then
	sram_write <= x"07DC0028";
end if;
if first_state_sram_input_id = 2774 then
	sram_write <= x"C05C0010";
end if;
if first_state_sram_input_id = 2775 then
	sram_write <= x"22440220";
end if;
if first_state_sram_input_id = 2776 then
	sram_write <= x"C07C0014";
end if;
if first_state_sram_input_id = 2777 then
	sram_write <= x"D4624000";
end if;
if first_state_sram_input_id = 2778 then
	sram_write <= x"82002B90";
end if;
if first_state_sram_input_id = 2779 then
	sram_write <= x"C03C0010";
end if;
if first_state_sram_input_id = 2780 then
	sram_write <= x"02220001";
end if;
if first_state_sram_input_id = 2781 then
	sram_write <= x"0240FFFF";
end if;
if first_state_sram_input_id = 2782 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2783 then
	sram_write <= x"03DC0028";
end if;
if first_state_sram_input_id = 2784 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2785 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2786 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 2787 then
	sram_write <= x"07DC0028";
end if;
if first_state_sram_input_id = 2788 then
	sram_write <= x"C05C0008";
end if;
if first_state_sram_input_id = 2789 then
	sram_write <= x"22440220";
end if;
if first_state_sram_input_id = 2790 then
	sram_write <= x"C07C000C";
end if;
if first_state_sram_input_id = 2791 then
	sram_write <= x"D4624000";
end if;
if first_state_sram_input_id = 2792 then
	sram_write <= x"82002BC8";
end if;
if first_state_sram_input_id = 2793 then
	sram_write <= x"C03C0008";
end if;
if first_state_sram_input_id = 2794 then
	sram_write <= x"02220001";
end if;
if first_state_sram_input_id = 2795 then
	sram_write <= x"0240FFFF";
end if;
if first_state_sram_input_id = 2796 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2797 then
	sram_write <= x"03DC0028";
end if;
if first_state_sram_input_id = 2798 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2799 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2800 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 2801 then
	sram_write <= x"07DC0028";
end if;
if first_state_sram_input_id = 2802 then
	sram_write <= x"C05C0000";
end if;
if first_state_sram_input_id = 2803 then
	sram_write <= x"22440220";
end if;
if first_state_sram_input_id = 2804 then
	sram_write <= x"C07C0004";
end if;
if first_state_sram_input_id = 2805 then
	sram_write <= x"D4624000";
end if;
if first_state_sram_input_id = 2806 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 2807 then
	sram_write <= x"C03C0000";
end if;
if first_state_sram_input_id = 2808 then
	sram_write <= x"02220001";
end if;
if first_state_sram_input_id = 2809 then
	sram_write <= x"0240FFFF";
end if;
if first_state_sram_input_id = 2810 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 2811 then
	sram_write <= x"C43C0000";
end if;
if first_state_sram_input_id = 2812 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2813 then
	sram_write <= x"03DC000C";
end if;
if first_state_sram_input_id = 2814 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2815 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2816 then
	sram_write <= x"82000794";
end if;
if first_state_sram_input_id = 2817 then
	sram_write <= x"07DC000C";
end if;
if first_state_sram_input_id = 2818 then
	sram_write <= x"0240FFFF";
end if;
if first_state_sram_input_id = 2819 then
	sram_write <= x"82242CE4";
end if;
if first_state_sram_input_id = 2820 then
	sram_write <= x"C43C0004";
end if;
if first_state_sram_input_id = 2821 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2822 then
	sram_write <= x"03DC0010";
end if;
if first_state_sram_input_id = 2823 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2824 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2825 then
	sram_write <= x"82000794";
end if;
if first_state_sram_input_id = 2826 then
	sram_write <= x"07DC0010";
end if;
if first_state_sram_input_id = 2827 then
	sram_write <= x"0240FFFF";
end if;
if first_state_sram_input_id = 2828 then
	sram_write <= x"82242CB4";
end if;
if first_state_sram_input_id = 2829 then
	sram_write <= x"C43C0008";
end if;
if first_state_sram_input_id = 2830 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2831 then
	sram_write <= x"03DC0014";
end if;
if first_state_sram_input_id = 2832 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2833 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2834 then
	sram_write <= x"82000794";
end if;
if first_state_sram_input_id = 2835 then
	sram_write <= x"07DC0014";
end if;
if first_state_sram_input_id = 2836 then
	sram_write <= x"0240FFFF";
end if;
if first_state_sram_input_id = 2837 then
	sram_write <= x"82242C88";
end if;
if first_state_sram_input_id = 2838 then
	sram_write <= x"02400003";
end if;
if first_state_sram_input_id = 2839 then
	sram_write <= x"C43C000C";
end if;
if first_state_sram_input_id = 2840 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2841 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 2842 then
	sram_write <= x"03DC0018";
end if;
if first_state_sram_input_id = 2843 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2844 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2845 then
	sram_write <= x"82002A44";
end if;
if first_state_sram_input_id = 2846 then
	sram_write <= x"07DC0018";
end if;
if first_state_sram_input_id = 2847 then
	sram_write <= x"C05C000C";
end if;
if first_state_sram_input_id = 2848 then
	sram_write <= x"C4420008";
end if;
if first_state_sram_input_id = 2849 then
	sram_write <= x"82002CA8";
end if;
if first_state_sram_input_id = 2850 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 2851 then
	sram_write <= x"0240FFFF";
end if;
if first_state_sram_input_id = 2852 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2853 then
	sram_write <= x"03DC0018";
end if;
if first_state_sram_input_id = 2854 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2855 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2856 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 2857 then
	sram_write <= x"07DC0018";
end if;
if first_state_sram_input_id = 2858 then
	sram_write <= x"C05C0008";
end if;
if first_state_sram_input_id = 2859 then
	sram_write <= x"C4420004";
end if;
if first_state_sram_input_id = 2860 then
	sram_write <= x"82002CD4";
end if;
if first_state_sram_input_id = 2861 then
	sram_write <= x"02200002";
end if;
if first_state_sram_input_id = 2862 then
	sram_write <= x"0240FFFF";
end if;
if first_state_sram_input_id = 2863 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2864 then
	sram_write <= x"03DC0018";
end if;
if first_state_sram_input_id = 2865 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2866 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2867 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 2868 then
	sram_write <= x"07DC0018";
end if;
if first_state_sram_input_id = 2869 then
	sram_write <= x"C05C0004";
end if;
if first_state_sram_input_id = 2870 then
	sram_write <= x"C4420000";
end if;
if first_state_sram_input_id = 2871 then
	sram_write <= x"00420000";
end if;
if first_state_sram_input_id = 2872 then
	sram_write <= x"82002D08";
end if;
if first_state_sram_input_id = 2873 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 2874 then
	sram_write <= x"0240FFFF";
end if;
if first_state_sram_input_id = 2875 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2876 then
	sram_write <= x"03DC0018";
end if;
if first_state_sram_input_id = 2877 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2878 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2879 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 2880 then
	sram_write <= x"07DC0018";
end if;
if first_state_sram_input_id = 2881 then
	sram_write <= x"00420000";
end if;
if first_state_sram_input_id = 2882 then
	sram_write <= x"C0240000";
end if;
if first_state_sram_input_id = 2883 then
	sram_write <= x"0260FFFF";
end if;
if first_state_sram_input_id = 2884 then
	sram_write <= x"82262E68";
end if;
if first_state_sram_input_id = 2885 then
	sram_write <= x"C03C0000";
end if;
if first_state_sram_input_id = 2886 then
	sram_write <= x"02620001";
end if;
if first_state_sram_input_id = 2887 then
	sram_write <= x"C45C0010";
end if;
if first_state_sram_input_id = 2888 then
	sram_write <= x"C47C0014";
end if;
if first_state_sram_input_id = 2889 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2890 then
	sram_write <= x"03DC0020";
end if;
if first_state_sram_input_id = 2891 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2892 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2893 then
	sram_write <= x"82000794";
end if;
if first_state_sram_input_id = 2894 then
	sram_write <= x"07DC0020";
end if;
if first_state_sram_input_id = 2895 then
	sram_write <= x"0240FFFF";
end if;
if first_state_sram_input_id = 2896 then
	sram_write <= x"82242DC8";
end if;
if first_state_sram_input_id = 2897 then
	sram_write <= x"C43C0018";
end if;
if first_state_sram_input_id = 2898 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2899 then
	sram_write <= x"03DC0024";
end if;
if first_state_sram_input_id = 2900 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2901 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2902 then
	sram_write <= x"82000794";
end if;
if first_state_sram_input_id = 2903 then
	sram_write <= x"07DC0024";
end if;
if first_state_sram_input_id = 2904 then
	sram_write <= x"0240FFFF";
end if;
if first_state_sram_input_id = 2905 then
	sram_write <= x"82242D98";
end if;
if first_state_sram_input_id = 2906 then
	sram_write <= x"02400002";
end if;
if first_state_sram_input_id = 2907 then
	sram_write <= x"C43C001C";
end if;
if first_state_sram_input_id = 2908 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2909 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 2910 then
	sram_write <= x"03DC0028";
end if;
if first_state_sram_input_id = 2911 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2912 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2913 then
	sram_write <= x"82002A44";
end if;
if first_state_sram_input_id = 2914 then
	sram_write <= x"07DC0028";
end if;
if first_state_sram_input_id = 2915 then
	sram_write <= x"C05C001C";
end if;
if first_state_sram_input_id = 2916 then
	sram_write <= x"C4420004";
end if;
if first_state_sram_input_id = 2917 then
	sram_write <= x"82002DB8";
end if;
if first_state_sram_input_id = 2918 then
	sram_write <= x"02200002";
end if;
if first_state_sram_input_id = 2919 then
	sram_write <= x"0240FFFF";
end if;
if first_state_sram_input_id = 2920 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2921 then
	sram_write <= x"03DC0028";
end if;
if first_state_sram_input_id = 2922 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2923 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2924 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 2925 then
	sram_write <= x"07DC0028";
end if;
if first_state_sram_input_id = 2926 then
	sram_write <= x"C05C0018";
end if;
if first_state_sram_input_id = 2927 then
	sram_write <= x"C4420000";
end if;
if first_state_sram_input_id = 2928 then
	sram_write <= x"00420000";
end if;
if first_state_sram_input_id = 2929 then
	sram_write <= x"82002DEC";
end if;
if first_state_sram_input_id = 2930 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 2931 then
	sram_write <= x"0240FFFF";
end if;
if first_state_sram_input_id = 2932 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2933 then
	sram_write <= x"03DC0028";
end if;
if first_state_sram_input_id = 2934 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2935 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2936 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 2937 then
	sram_write <= x"07DC0028";
end if;
if first_state_sram_input_id = 2938 then
	sram_write <= x"00420000";
end if;
if first_state_sram_input_id = 2939 then
	sram_write <= x"C0240000";
end if;
if first_state_sram_input_id = 2940 then
	sram_write <= x"0260FFFF";
end if;
if first_state_sram_input_id = 2941 then
	sram_write <= x"82262E34";
end if;
if first_state_sram_input_id = 2942 then
	sram_write <= x"C03C0014";
end if;
if first_state_sram_input_id = 2943 then
	sram_write <= x"02620001";
end if;
if first_state_sram_input_id = 2944 then
	sram_write <= x"C45C0020";
end if;
if first_state_sram_input_id = 2945 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2946 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 2947 then
	sram_write <= x"03DC002C";
end if;
if first_state_sram_input_id = 2948 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2949 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2950 then
	sram_write <= x"82002BEC";
end if;
if first_state_sram_input_id = 2951 then
	sram_write <= x"07DC002C";
end if;
if first_state_sram_input_id = 2952 then
	sram_write <= x"C05C0014";
end if;
if first_state_sram_input_id = 2953 then
	sram_write <= x"22440220";
end if;
if first_state_sram_input_id = 2954 then
	sram_write <= x"C07C0020";
end if;
if first_state_sram_input_id = 2955 then
	sram_write <= x"D4624000";
end if;
if first_state_sram_input_id = 2956 then
	sram_write <= x"82002E54";
end if;
if first_state_sram_input_id = 2957 then
	sram_write <= x"C03C0014";
end if;
if first_state_sram_input_id = 2958 then
	sram_write <= x"02220001";
end if;
if first_state_sram_input_id = 2959 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2960 then
	sram_write <= x"03DC002C";
end if;
if first_state_sram_input_id = 2961 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2962 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2963 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 2964 then
	sram_write <= x"07DC002C";
end if;
if first_state_sram_input_id = 2965 then
	sram_write <= x"C05C0000";
end if;
if first_state_sram_input_id = 2966 then
	sram_write <= x"22440220";
end if;
if first_state_sram_input_id = 2967 then
	sram_write <= x"C07C0010";
end if;
if first_state_sram_input_id = 2968 then
	sram_write <= x"D4624000";
end if;
if first_state_sram_input_id = 2969 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 2970 then
	sram_write <= x"C03C0000";
end if;
if first_state_sram_input_id = 2971 then
	sram_write <= x"02220001";
end if;
if first_state_sram_input_id = 2972 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 2973 then
	sram_write <= x"C43C0000";
end if;
if first_state_sram_input_id = 2974 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2975 then
	sram_write <= x"03DC000C";
end if;
if first_state_sram_input_id = 2976 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2977 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2978 then
	sram_write <= x"82000794";
end if;
if first_state_sram_input_id = 2979 then
	sram_write <= x"07DC000C";
end if;
if first_state_sram_input_id = 2980 then
	sram_write <= x"0240FFFF";
end if;
if first_state_sram_input_id = 2981 then
	sram_write <= x"82242F68";
end if;
if first_state_sram_input_id = 2982 then
	sram_write <= x"C43C0004";
end if;
if first_state_sram_input_id = 2983 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2984 then
	sram_write <= x"03DC0010";
end if;
if first_state_sram_input_id = 2985 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2986 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2987 then
	sram_write <= x"82000794";
end if;
if first_state_sram_input_id = 2988 then
	sram_write <= x"07DC0010";
end if;
if first_state_sram_input_id = 2989 then
	sram_write <= x"0240FFFF";
end if;
if first_state_sram_input_id = 2990 then
	sram_write <= x"82242F3C";
end if;
if first_state_sram_input_id = 2991 then
	sram_write <= x"C43C0008";
end if;
if first_state_sram_input_id = 2992 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 2993 then
	sram_write <= x"03DC0014";
end if;
if first_state_sram_input_id = 2994 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 2995 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 2996 then
	sram_write <= x"82000794";
end if;
if first_state_sram_input_id = 2997 then
	sram_write <= x"07DC0014";
end if;
if first_state_sram_input_id = 2998 then
	sram_write <= x"0240FFFF";
end if;
if first_state_sram_input_id = 2999 then
	sram_write <= x"82242F10";
end if;
if first_state_sram_input_id = 3000 then
	sram_write <= x"02400003";
end if;
if first_state_sram_input_id = 3001 then
	sram_write <= x"C43C000C";
end if;
if first_state_sram_input_id = 3002 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 3003 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 3004 then
	sram_write <= x"03DC0018";
end if;
if first_state_sram_input_id = 3005 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 3006 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 3007 then
	sram_write <= x"82002A44";
end if;
if first_state_sram_input_id = 3008 then
	sram_write <= x"07DC0018";
end if;
if first_state_sram_input_id = 3009 then
	sram_write <= x"C05C000C";
end if;
if first_state_sram_input_id = 3010 then
	sram_write <= x"C4420008";
end if;
if first_state_sram_input_id = 3011 then
	sram_write <= x"82002F30";
end if;
if first_state_sram_input_id = 3012 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 3013 then
	sram_write <= x"0240FFFF";
end if;
if first_state_sram_input_id = 3014 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 3015 then
	sram_write <= x"03DC0018";
end if;
if first_state_sram_input_id = 3016 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 3017 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 3018 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 3019 then
	sram_write <= x"07DC0018";
end if;
if first_state_sram_input_id = 3020 then
	sram_write <= x"C05C0008";
end if;
if first_state_sram_input_id = 3021 then
	sram_write <= x"C4420004";
end if;
if first_state_sram_input_id = 3022 then
	sram_write <= x"82002F5C";
end if;
if first_state_sram_input_id = 3023 then
	sram_write <= x"02200002";
end if;
if first_state_sram_input_id = 3024 then
	sram_write <= x"0240FFFF";
end if;
if first_state_sram_input_id = 3025 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 3026 then
	sram_write <= x"03DC0018";
end if;
if first_state_sram_input_id = 3027 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 3028 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 3029 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 3030 then
	sram_write <= x"07DC0018";
end if;
if first_state_sram_input_id = 3031 then
	sram_write <= x"C05C0004";
end if;
if first_state_sram_input_id = 3032 then
	sram_write <= x"C4420000";
end if;
if first_state_sram_input_id = 3033 then
	sram_write <= x"82002F88";
end if;
if first_state_sram_input_id = 3034 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 3035 then
	sram_write <= x"0240FFFF";
end if;
if first_state_sram_input_id = 3036 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 3037 then
	sram_write <= x"03DC0018";
end if;
if first_state_sram_input_id = 3038 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 3039 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 3040 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 3041 then
	sram_write <= x"07DC0018";
end if;
if first_state_sram_input_id = 3042 then
	sram_write <= x"C0420000";
end if;
if first_state_sram_input_id = 3043 then
	sram_write <= x"0260FFFF";
end if;
if first_state_sram_input_id = 3044 then
	sram_write <= x"82463178";
end if;
if first_state_sram_input_id = 3045 then
	sram_write <= x"024001E0";
end if;
if first_state_sram_input_id = 3046 then
	sram_write <= x"C07C0000";
end if;
if first_state_sram_input_id = 3047 then
	sram_write <= x"22860220";
end if;
if first_state_sram_input_id = 3048 then
	sram_write <= x"D4248000";
end if;
if first_state_sram_input_id = 3049 then
	sram_write <= x"02260001";
end if;
if first_state_sram_input_id = 3050 then
	sram_write <= x"C45C0010";
end if;
if first_state_sram_input_id = 3051 then
	sram_write <= x"C43C0014";
end if;
if first_state_sram_input_id = 3052 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 3053 then
	sram_write <= x"03DC0020";
end if;
if first_state_sram_input_id = 3054 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 3055 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 3056 then
	sram_write <= x"82000794";
end if;
if first_state_sram_input_id = 3057 then
	sram_write <= x"07DC0020";
end if;
if first_state_sram_input_id = 3058 then
	sram_write <= x"0240FFFF";
end if;
if first_state_sram_input_id = 3059 then
	sram_write <= x"82243050";
end if;
if first_state_sram_input_id = 3060 then
	sram_write <= x"C43C0018";
end if;
if first_state_sram_input_id = 3061 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 3062 then
	sram_write <= x"03DC0024";
end if;
if first_state_sram_input_id = 3063 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 3064 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 3065 then
	sram_write <= x"82000794";
end if;
if first_state_sram_input_id = 3066 then
	sram_write <= x"07DC0024";
end if;
if first_state_sram_input_id = 3067 then
	sram_write <= x"0240FFFF";
end if;
if first_state_sram_input_id = 3068 then
	sram_write <= x"82243024";
end if;
if first_state_sram_input_id = 3069 then
	sram_write <= x"02400002";
end if;
if first_state_sram_input_id = 3070 then
	sram_write <= x"C43C001C";
end if;
if first_state_sram_input_id = 3071 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 3072 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 3073 then
	sram_write <= x"03DC0028";
end if;
if first_state_sram_input_id = 3074 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 3075 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 3076 then
	sram_write <= x"82002A44";
end if;
if first_state_sram_input_id = 3077 then
	sram_write <= x"07DC0028";
end if;
if first_state_sram_input_id = 3078 then
	sram_write <= x"C05C001C";
end if;
if first_state_sram_input_id = 3079 then
	sram_write <= x"C4420004";
end if;
if first_state_sram_input_id = 3080 then
	sram_write <= x"82003044";
end if;
if first_state_sram_input_id = 3081 then
	sram_write <= x"02200002";
end if;
if first_state_sram_input_id = 3082 then
	sram_write <= x"0240FFFF";
end if;
if first_state_sram_input_id = 3083 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 3084 then
	sram_write <= x"03DC0028";
end if;
if first_state_sram_input_id = 3085 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 3086 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 3087 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 3088 then
	sram_write <= x"07DC0028";
end if;
if first_state_sram_input_id = 3089 then
	sram_write <= x"C05C0018";
end if;
if first_state_sram_input_id = 3090 then
	sram_write <= x"C4420000";
end if;
if first_state_sram_input_id = 3091 then
	sram_write <= x"82003070";
end if;
if first_state_sram_input_id = 3092 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 3093 then
	sram_write <= x"0240FFFF";
end if;
if first_state_sram_input_id = 3094 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 3095 then
	sram_write <= x"03DC0028";
end if;
if first_state_sram_input_id = 3096 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 3097 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 3098 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 3099 then
	sram_write <= x"07DC0028";
end if;
if first_state_sram_input_id = 3100 then
	sram_write <= x"C0420000";
end if;
if first_state_sram_input_id = 3101 then
	sram_write <= x"0260FFFF";
end if;
if first_state_sram_input_id = 3102 then
	sram_write <= x"82463174";
end if;
if first_state_sram_input_id = 3103 then
	sram_write <= x"C05C0014";
end if;
if first_state_sram_input_id = 3104 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 3105 then
	sram_write <= x"C09C0010";
end if;
if first_state_sram_input_id = 3106 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 3107 then
	sram_write <= x"02240001";
end if;
if first_state_sram_input_id = 3108 then
	sram_write <= x"C43C0020";
end if;
if first_state_sram_input_id = 3109 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 3110 then
	sram_write <= x"03DC002C";
end if;
if first_state_sram_input_id = 3111 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 3112 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 3113 then
	sram_write <= x"82000794";
end if;
if first_state_sram_input_id = 3114 then
	sram_write <= x"07DC002C";
end if;
if first_state_sram_input_id = 3115 then
	sram_write <= x"0240FFFF";
end if;
if first_state_sram_input_id = 3116 then
	sram_write <= x"822430E4";
end if;
if first_state_sram_input_id = 3117 then
	sram_write <= x"02400001";
end if;
if first_state_sram_input_id = 3118 then
	sram_write <= x"C43C0024";
end if;
if first_state_sram_input_id = 3119 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 3120 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 3121 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 3122 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 3123 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 3124 then
	sram_write <= x"82002A44";
end if;
if first_state_sram_input_id = 3125 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 3126 then
	sram_write <= x"C05C0024";
end if;
if first_state_sram_input_id = 3127 then
	sram_write <= x"C4420000";
end if;
if first_state_sram_input_id = 3128 then
	sram_write <= x"82003104";
end if;
if first_state_sram_input_id = 3129 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 3130 then
	sram_write <= x"0240FFFF";
end if;
if first_state_sram_input_id = 3131 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 3132 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 3133 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 3134 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 3135 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 3136 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 3137 then
	sram_write <= x"C0420000";
end if;
if first_state_sram_input_id = 3138 then
	sram_write <= x"0260FFFF";
end if;
if first_state_sram_input_id = 3139 then
	sram_write <= x"82463170";
end if;
if first_state_sram_input_id = 3140 then
	sram_write <= x"C05C0020";
end if;
if first_state_sram_input_id = 3141 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 3142 then
	sram_write <= x"C09C0010";
end if;
if first_state_sram_input_id = 3143 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 3144 then
	sram_write <= x"02240001";
end if;
if first_state_sram_input_id = 3145 then
	sram_write <= x"02400000";
end if;
if first_state_sram_input_id = 3146 then
	sram_write <= x"C43C0028";
end if;
if first_state_sram_input_id = 3147 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 3148 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 3149 then
	sram_write <= x"03DC0034";
end if;
if first_state_sram_input_id = 3150 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 3151 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 3152 then
	sram_write <= x"82002A44";
end if;
if first_state_sram_input_id = 3153 then
	sram_write <= x"07DC0034";
end if;
if first_state_sram_input_id = 3154 then
	sram_write <= x"C0420000";
end if;
if first_state_sram_input_id = 3155 then
	sram_write <= x"0260FFFF";
end if;
if first_state_sram_input_id = 3156 then
	sram_write <= x"8246316C";
end if;
if first_state_sram_input_id = 3157 then
	sram_write <= x"C05C0028";
end if;
if first_state_sram_input_id = 3158 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 3159 then
	sram_write <= x"C09C0010";
end if;
if first_state_sram_input_id = 3160 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 3161 then
	sram_write <= x"02240001";
end if;
if first_state_sram_input_id = 3162 then
	sram_write <= x"82002E74";
end if;
if first_state_sram_input_id = 3163 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 3164 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 3165 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 3166 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 3167 then
	sram_write <= x"22C60220";
end if;
if first_state_sram_input_id = 3168 then
	sram_write <= x"D884C000";
end if;
if first_state_sram_input_id = 3169 then
	sram_write <= x"8A80329C";
end if;
if first_state_sram_input_id = 3170 then
	sram_write <= x"C0C20010";
end if;
if first_state_sram_input_id = 3171 then
	sram_write <= x"C0220018";
end if;
if first_state_sram_input_id = 3172 then
	sram_write <= x"8E80319C";
end if;
if first_state_sram_input_id = 3173 then
	sram_write <= x"02E00000";
end if;
if first_state_sram_input_id = 3174 then
	sram_write <= x"820031A0";
end if;
if first_state_sram_input_id = 3175 then
	sram_write <= x"02E00001";
end if;
if first_state_sram_input_id = 3176 then
	sram_write <= x"822031B8";
end if;
if first_state_sram_input_id = 3177 then
	sram_write <= x"8E8031B0";
end if;
if first_state_sram_input_id = 3178 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 3179 then
	sram_write <= x"820031B4";
end if;
if first_state_sram_input_id = 3180 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 3181 then
	sram_write <= x"820031BC";
end if;
if first_state_sram_input_id = 3182 then
	sram_write <= x"002E0000";
end if;
if first_state_sram_input_id = 3183 then
	sram_write <= x"22660220";
end if;
if first_state_sram_input_id = 3184 then
	sram_write <= x"D8AC6000";
end if;
if first_state_sram_input_id = 3185 then
	sram_write <= x"822031CC";
end if;
if first_state_sram_input_id = 3186 then
	sram_write <= x"820031D0";
end if;
if first_state_sram_input_id = 3187 then
	sram_write <= x"44A0A000";
end if;
if first_state_sram_input_id = 3188 then
	sram_write <= x"442A2000";
end if;
if first_state_sram_input_id = 3189 then
	sram_write <= x"CC7C0000";
end if;
if first_state_sram_input_id = 3190 then
	sram_write <= x"C4BC0008";
end if;
if first_state_sram_input_id = 3191 then
	sram_write <= x"C4DC000C";
end if;
if first_state_sram_input_id = 3192 then
	sram_write <= x"CC5C0010";
end if;
if first_state_sram_input_id = 3193 then
	sram_write <= x"C45C0018";
end if;
if first_state_sram_input_id = 3194 then
	sram_write <= x"C49C001C";
end if;
if first_state_sram_input_id = 3195 then
	sram_write <= x"CC3C0020";
end if;
if first_state_sram_input_id = 3196 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 3197 then
	sram_write <= x"40208000";
end if;
if first_state_sram_input_id = 3198 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 3199 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 3200 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 3201 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 3202 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 3203 then
	sram_write <= x"C85C0020";
end if;
if first_state_sram_input_id = 3204 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 3205 then
	sram_write <= x"C03C001C";
end if;
if first_state_sram_input_id = 3206 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 3207 then
	sram_write <= x"C07C0018";
end if;
if first_state_sram_input_id = 3208 then
	sram_write <= x"D8464000";
end if;
if first_state_sram_input_id = 3209 then
	sram_write <= x"48424000";
end if;
if first_state_sram_input_id = 3210 then
	sram_write <= x"C87C0010";
end if;
if first_state_sram_input_id = 3211 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 3212 then
	sram_write <= x"8E403238";
end if;
if first_state_sram_input_id = 3213 then
	sram_write <= x"8200323C";
end if;
if first_state_sram_input_id = 3214 then
	sram_write <= x"44404000";
end if;
if first_state_sram_input_id = 3215 then
	sram_write <= x"22220220";
end if;
if first_state_sram_input_id = 3216 then
	sram_write <= x"C05C000C";
end if;
if first_state_sram_input_id = 3217 then
	sram_write <= x"D8642000";
end if;
if first_state_sram_input_id = 3218 then
	sram_write <= x"8E463254";
end if;
if first_state_sram_input_id = 3219 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 3220 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 3221 then
	sram_write <= x"C03C0008";
end if;
if first_state_sram_input_id = 3222 then
	sram_write <= x"22820220";
end if;
if first_state_sram_input_id = 3223 then
	sram_write <= x"D8468000";
end if;
if first_state_sram_input_id = 3224 then
	sram_write <= x"48424000";
end if;
if first_state_sram_input_id = 3225 then
	sram_write <= x"C87C0000";
end if;
if first_state_sram_input_id = 3226 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 3227 then
	sram_write <= x"8E403274";
end if;
if first_state_sram_input_id = 3228 then
	sram_write <= x"82003278";
end if;
if first_state_sram_input_id = 3229 then
	sram_write <= x"44404000";
end if;
if first_state_sram_input_id = 3230 then
	sram_write <= x"22220220";
end if;
if first_state_sram_input_id = 3231 then
	sram_write <= x"D8642000";
end if;
if first_state_sram_input_id = 3232 then
	sram_write <= x"8E46328C";
end if;
if first_state_sram_input_id = 3233 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 3234 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 3235 then
	sram_write <= x"022002AC";
end if;
if first_state_sram_input_id = 3236 then
	sram_write <= x"CC220000";
end if;
if first_state_sram_input_id = 3237 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 3238 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 3239 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 3240 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 3241 then
	sram_write <= x"C0220010";
end if;
if first_state_sram_input_id = 3242 then
	sram_write <= x"C8840000";
end if;
if first_state_sram_input_id = 3243 then
	sram_write <= x"C8A20000";
end if;
if first_state_sram_input_id = 3244 then
	sram_write <= x"4888A000";
end if;
if first_state_sram_input_id = 3245 then
	sram_write <= x"C8A40004";
end if;
if first_state_sram_input_id = 3246 then
	sram_write <= x"C8C20004";
end if;
if first_state_sram_input_id = 3247 then
	sram_write <= x"48AAC000";
end if;
if first_state_sram_input_id = 3248 then
	sram_write <= x"4088A000";
end if;
if first_state_sram_input_id = 3249 then
	sram_write <= x"C8A40008";
end if;
if first_state_sram_input_id = 3250 then
	sram_write <= x"C8C20008";
end if;
if first_state_sram_input_id = 3251 then
	sram_write <= x"48AAC000";
end if;
if first_state_sram_input_id = 3252 then
	sram_write <= x"4088A000";
end if;
if first_state_sram_input_id = 3253 then
	sram_write <= x"8E0832E0";
end if;
if first_state_sram_input_id = 3254 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 3255 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 3256 then
	sram_write <= x"024002AC";
end if;
if first_state_sram_input_id = 3257 then
	sram_write <= x"C8A20000";
end if;
if first_state_sram_input_id = 3258 then
	sram_write <= x"482A2000";
end if;
if first_state_sram_input_id = 3259 then
	sram_write <= x"C8A20004";
end if;
if first_state_sram_input_id = 3260 then
	sram_write <= x"484A4000";
end if;
if first_state_sram_input_id = 3261 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 3262 then
	sram_write <= x"C8420008";
end if;
if first_state_sram_input_id = 3263 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 3264 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 3265 then
	sram_write <= x"44202000";
end if;
if first_state_sram_input_id = 3266 then
	sram_write <= x"C45C0000";
end if;
if first_state_sram_input_id = 3267 then
	sram_write <= x"CC3C0008";
end if;
if first_state_sram_input_id = 3268 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 3269 then
	sram_write <= x"40208000";
end if;
if first_state_sram_input_id = 3270 then
	sram_write <= x"03DC0018";
end if;
if first_state_sram_input_id = 3271 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 3272 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 3273 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 3274 then
	sram_write <= x"07DC0018";
end if;
if first_state_sram_input_id = 3275 then
	sram_write <= x"C85C0008";
end if;
if first_state_sram_input_id = 3276 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 3277 then
	sram_write <= x"C03C0000";
end if;
if first_state_sram_input_id = 3278 then
	sram_write <= x"CC220000";
end if;
if first_state_sram_input_id = 3279 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 3280 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 3281 then
	sram_write <= x"48822000";
end if;
if first_state_sram_input_id = 3282 then
	sram_write <= x"C0420010";
end if;
if first_state_sram_input_id = 3283 then
	sram_write <= x"C8A40000";
end if;
if first_state_sram_input_id = 3284 then
	sram_write <= x"4888A000";
end if;
if first_state_sram_input_id = 3285 then
	sram_write <= x"48A44000";
end if;
if first_state_sram_input_id = 3286 then
	sram_write <= x"C0420010";
end if;
if first_state_sram_input_id = 3287 then
	sram_write <= x"C8C40004";
end if;
if first_state_sram_input_id = 3288 then
	sram_write <= x"48AAC000";
end if;
if first_state_sram_input_id = 3289 then
	sram_write <= x"4088A000";
end if;
if first_state_sram_input_id = 3290 then
	sram_write <= x"48A66000";
end if;
if first_state_sram_input_id = 3291 then
	sram_write <= x"C0420010";
end if;
if first_state_sram_input_id = 3292 then
	sram_write <= x"C8C40008";
end if;
if first_state_sram_input_id = 3293 then
	sram_write <= x"48AAC000";
end if;
if first_state_sram_input_id = 3294 then
	sram_write <= x"4088A000";
end if;
if first_state_sram_input_id = 3295 then
	sram_write <= x"C042000C";
end if;
if first_state_sram_input_id = 3296 then
	sram_write <= x"824033C4";
end if;
if first_state_sram_input_id = 3297 then
	sram_write <= x"48A46000";
end if;
if first_state_sram_input_id = 3298 then
	sram_write <= x"C0420024";
end if;
if first_state_sram_input_id = 3299 then
	sram_write <= x"C8C40000";
end if;
if first_state_sram_input_id = 3300 then
	sram_write <= x"48AAC000";
end if;
if first_state_sram_input_id = 3301 then
	sram_write <= x"4088A000";
end if;
if first_state_sram_input_id = 3302 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 3303 then
	sram_write <= x"C0420024";
end if;
if first_state_sram_input_id = 3304 then
	sram_write <= x"C8A40004";
end if;
if first_state_sram_input_id = 3305 then
	sram_write <= x"4866A000";
end if;
if first_state_sram_input_id = 3306 then
	sram_write <= x"40686000";
end if;
if first_state_sram_input_id = 3307 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 3308 then
	sram_write <= x"C0220024";
end if;
if first_state_sram_input_id = 3309 then
	sram_write <= x"C8420008";
end if;
if first_state_sram_input_id = 3310 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 3311 then
	sram_write <= x"40262000";
end if;
if first_state_sram_input_id = 3312 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 3313 then
	sram_write <= x"40208000";
end if;
if first_state_sram_input_id = 3314 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 3315 then
	sram_write <= x"48E28000";
end if;
if first_state_sram_input_id = 3316 then
	sram_write <= x"C0420010";
end if;
if first_state_sram_input_id = 3317 then
	sram_write <= x"C9040000";
end if;
if first_state_sram_input_id = 3318 then
	sram_write <= x"48EF0000";
end if;
if first_state_sram_input_id = 3319 then
	sram_write <= x"4904A000";
end if;
if first_state_sram_input_id = 3320 then
	sram_write <= x"C0420010";
end if;
if first_state_sram_input_id = 3321 then
	sram_write <= x"C9240004";
end if;
if first_state_sram_input_id = 3322 then
	sram_write <= x"49112000";
end if;
if first_state_sram_input_id = 3323 then
	sram_write <= x"40EF0000";
end if;
if first_state_sram_input_id = 3324 then
	sram_write <= x"4906C000";
end if;
if first_state_sram_input_id = 3325 then
	sram_write <= x"C0420010";
end if;
if first_state_sram_input_id = 3326 then
	sram_write <= x"C9240008";
end if;
if first_state_sram_input_id = 3327 then
	sram_write <= x"49112000";
end if;
if first_state_sram_input_id = 3328 then
	sram_write <= x"40EF0000";
end if;
if first_state_sram_input_id = 3329 then
	sram_write <= x"C042000C";
end if;
if first_state_sram_input_id = 3330 then
	sram_write <= x"82403498";
end if;
if first_state_sram_input_id = 3331 then
	sram_write <= x"4906A000";
end if;
if first_state_sram_input_id = 3332 then
	sram_write <= x"4924C000";
end if;
if first_state_sram_input_id = 3333 then
	sram_write <= x"41112000";
end if;
if first_state_sram_input_id = 3334 then
	sram_write <= x"C0420024";
end if;
if first_state_sram_input_id = 3335 then
	sram_write <= x"C9240000";
end if;
if first_state_sram_input_id = 3336 then
	sram_write <= x"49112000";
end if;
if first_state_sram_input_id = 3337 then
	sram_write <= x"48C2C000";
end if;
if first_state_sram_input_id = 3338 then
	sram_write <= x"48668000";
end if;
if first_state_sram_input_id = 3339 then
	sram_write <= x"406C6000";
end if;
if first_state_sram_input_id = 3340 then
	sram_write <= x"C0420024";
end if;
if first_state_sram_input_id = 3341 then
	sram_write <= x"C8C40004";
end if;
if first_state_sram_input_id = 3342 then
	sram_write <= x"4866C000";
end if;
if first_state_sram_input_id = 3343 then
	sram_write <= x"40706000";
end if;
if first_state_sram_input_id = 3344 then
	sram_write <= x"4822A000";
end if;
if first_state_sram_input_id = 3345 then
	sram_write <= x"48448000";
end if;
if first_state_sram_input_id = 3346 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 3347 then
	sram_write <= x"C0220024";
end if;
if first_state_sram_input_id = 3348 then
	sram_write <= x"C8420008";
end if;
if first_state_sram_input_id = 3349 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 3350 then
	sram_write <= x"40262000";
end if;
if first_state_sram_input_id = 3351 then
	sram_write <= x"C8400080";
end if;
if first_state_sram_input_id = 3352 then
	sram_write <= x"CCFC0000";
end if;
if first_state_sram_input_id = 3353 then
	sram_write <= x"CC3C0008";
end if;
if first_state_sram_input_id = 3354 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 3355 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 3356 then
	sram_write <= x"03DC0018";
end if;
if first_state_sram_input_id = 3357 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 3358 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 3359 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 3360 then
	sram_write <= x"07DC0018";
end if;
if first_state_sram_input_id = 3361 then
	sram_write <= x"C85C0008";
end if;
if first_state_sram_input_id = 3362 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 3363 then
	sram_write <= x"C85C0000";
end if;
if first_state_sram_input_id = 3364 then
	sram_write <= x"40242000";
end if;
if first_state_sram_input_id = 3365 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 3366 then
	sram_write <= x"4020E000";
end if;
if first_state_sram_input_id = 3367 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 3368 then
	sram_write <= x"C8840000";
end if;
if first_state_sram_input_id = 3369 then
	sram_write <= x"C8A40004";
end if;
if first_state_sram_input_id = 3370 then
	sram_write <= x"C8C40008";
end if;
if first_state_sram_input_id = 3371 then
	sram_write <= x"48E88000";
end if;
if first_state_sram_input_id = 3372 then
	sram_write <= x"C0620010";
end if;
if first_state_sram_input_id = 3373 then
	sram_write <= x"C9060000";
end if;
if first_state_sram_input_id = 3374 then
	sram_write <= x"48EF0000";
end if;
if first_state_sram_input_id = 3375 then
	sram_write <= x"490AA000";
end if;
if first_state_sram_input_id = 3376 then
	sram_write <= x"C0620010";
end if;
if first_state_sram_input_id = 3377 then
	sram_write <= x"C9260004";
end if;
if first_state_sram_input_id = 3378 then
	sram_write <= x"49112000";
end if;
if first_state_sram_input_id = 3379 then
	sram_write <= x"40EF0000";
end if;
if first_state_sram_input_id = 3380 then
	sram_write <= x"490CC000";
end if;
if first_state_sram_input_id = 3381 then
	sram_write <= x"C0620010";
end if;
if first_state_sram_input_id = 3382 then
	sram_write <= x"C9260008";
end if;
if first_state_sram_input_id = 3383 then
	sram_write <= x"49112000";
end if;
if first_state_sram_input_id = 3384 then
	sram_write <= x"40EF0000";
end if;
if first_state_sram_input_id = 3385 then
	sram_write <= x"C062000C";
end if;
if first_state_sram_input_id = 3386 then
	sram_write <= x"8260352C";
end if;
if first_state_sram_input_id = 3387 then
	sram_write <= x"490AC000";
end if;
if first_state_sram_input_id = 3388 then
	sram_write <= x"C0620024";
end if;
if first_state_sram_input_id = 3389 then
	sram_write <= x"C9260000";
end if;
if first_state_sram_input_id = 3390 then
	sram_write <= x"49112000";
end if;
if first_state_sram_input_id = 3391 then
	sram_write <= x"40EF0000";
end if;
if first_state_sram_input_id = 3392 then
	sram_write <= x"48CC8000";
end if;
if first_state_sram_input_id = 3393 then
	sram_write <= x"C0620024";
end if;
if first_state_sram_input_id = 3394 then
	sram_write <= x"C9060004";
end if;
if first_state_sram_input_id = 3395 then
	sram_write <= x"48CD0000";
end if;
if first_state_sram_input_id = 3396 then
	sram_write <= x"40CEC000";
end if;
if first_state_sram_input_id = 3397 then
	sram_write <= x"4888A000";
end if;
if first_state_sram_input_id = 3398 then
	sram_write <= x"C0620024";
end if;
if first_state_sram_input_id = 3399 then
	sram_write <= x"C8A60008";
end if;
if first_state_sram_input_id = 3400 then
	sram_write <= x"4888A000";
end if;
if first_state_sram_input_id = 3401 then
	sram_write <= x"408C8000";
end if;
if first_state_sram_input_id = 3402 then
	sram_write <= x"82003530";
end if;
if first_state_sram_input_id = 3403 then
	sram_write <= x"4080E000";
end if;
if first_state_sram_input_id = 3404 then
	sram_write <= x"8A8036CC";
end if;
if first_state_sram_input_id = 3405 then
	sram_write <= x"C8A40000";
end if;
if first_state_sram_input_id = 3406 then
	sram_write <= x"C8C40004";
end if;
if first_state_sram_input_id = 3407 then
	sram_write <= x"C8E40008";
end if;
if first_state_sram_input_id = 3408 then
	sram_write <= x"CC9C0000";
end if;
if first_state_sram_input_id = 3409 then
	sram_write <= x"CC7C0008";
end if;
if first_state_sram_input_id = 3410 then
	sram_write <= x"CC5C0010";
end if;
if first_state_sram_input_id = 3411 then
	sram_write <= x"C43C0018";
end if;
if first_state_sram_input_id = 3412 then
	sram_write <= x"CC3C0020";
end if;
if first_state_sram_input_id = 3413 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 3414 then
	sram_write <= x"40802000";
end if;
if first_state_sram_input_id = 3415 then
	sram_write <= x"4020A000";
end if;
if first_state_sram_input_id = 3416 then
	sram_write <= x"40A04000";
end if;
if first_state_sram_input_id = 3417 then
	sram_write <= x"4040C000";
end if;
if first_state_sram_input_id = 3418 then
	sram_write <= x"40C06000";
end if;
if first_state_sram_input_id = 3419 then
	sram_write <= x"4060E000";
end if;
if first_state_sram_input_id = 3420 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 3421 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 3422 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 3423 then
	sram_write <= x"820033CC";
end if;
if first_state_sram_input_id = 3424 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 3425 then
	sram_write <= x"C85C0020";
end if;
if first_state_sram_input_id = 3426 then
	sram_write <= x"48644000";
end if;
if first_state_sram_input_id = 3427 then
	sram_write <= x"C03C0018";
end if;
if first_state_sram_input_id = 3428 then
	sram_write <= x"C0420010";
end if;
if first_state_sram_input_id = 3429 then
	sram_write <= x"C8840000";
end if;
if first_state_sram_input_id = 3430 then
	sram_write <= x"48668000";
end if;
if first_state_sram_input_id = 3431 then
	sram_write <= x"C89C0010";
end if;
if first_state_sram_input_id = 3432 then
	sram_write <= x"48A88000";
end if;
if first_state_sram_input_id = 3433 then
	sram_write <= x"C0420010";
end if;
if first_state_sram_input_id = 3434 then
	sram_write <= x"C8C40004";
end if;
if first_state_sram_input_id = 3435 then
	sram_write <= x"48AAC000";
end if;
if first_state_sram_input_id = 3436 then
	sram_write <= x"4066A000";
end if;
if first_state_sram_input_id = 3437 then
	sram_write <= x"C8BC0008";
end if;
if first_state_sram_input_id = 3438 then
	sram_write <= x"48CAA000";
end if;
if first_state_sram_input_id = 3439 then
	sram_write <= x"C0420010";
end if;
if first_state_sram_input_id = 3440 then
	sram_write <= x"C8E40008";
end if;
if first_state_sram_input_id = 3441 then
	sram_write <= x"48CCE000";
end if;
if first_state_sram_input_id = 3442 then
	sram_write <= x"4066C000";
end if;
if first_state_sram_input_id = 3443 then
	sram_write <= x"C042000C";
end if;
if first_state_sram_input_id = 3444 then
	sram_write <= x"82403614";
end if;
if first_state_sram_input_id = 3445 then
	sram_write <= x"48C8A000";
end if;
if first_state_sram_input_id = 3446 then
	sram_write <= x"C0420024";
end if;
if first_state_sram_input_id = 3447 then
	sram_write <= x"C8E40000";
end if;
if first_state_sram_input_id = 3448 then
	sram_write <= x"48CCE000";
end if;
if first_state_sram_input_id = 3449 then
	sram_write <= x"4066C000";
end if;
if first_state_sram_input_id = 3450 then
	sram_write <= x"48AA4000";
end if;
if first_state_sram_input_id = 3451 then
	sram_write <= x"C0420024";
end if;
if first_state_sram_input_id = 3452 then
	sram_write <= x"C8C40004";
end if;
if first_state_sram_input_id = 3453 then
	sram_write <= x"48AAC000";
end if;
if first_state_sram_input_id = 3454 then
	sram_write <= x"4066A000";
end if;
if first_state_sram_input_id = 3455 then
	sram_write <= x"48448000";
end if;
if first_state_sram_input_id = 3456 then
	sram_write <= x"C0420024";
end if;
if first_state_sram_input_id = 3457 then
	sram_write <= x"C8840008";
end if;
if first_state_sram_input_id = 3458 then
	sram_write <= x"48448000";
end if;
if first_state_sram_input_id = 3459 then
	sram_write <= x"40464000";
end if;
if first_state_sram_input_id = 3460 then
	sram_write <= x"82003618";
end if;
if first_state_sram_input_id = 3461 then
	sram_write <= x"40406000";
end if;
if first_state_sram_input_id = 3462 then
	sram_write <= x"C0420004";
end if;
if first_state_sram_input_id = 3463 then
	sram_write <= x"02600003";
end if;
if first_state_sram_input_id = 3464 then
	sram_write <= x"82463628";
end if;
if first_state_sram_input_id = 3465 then
	sram_write <= x"82003630";
end if;
if first_state_sram_input_id = 3466 then
	sram_write <= x"C86000A8";
end if;
if first_state_sram_input_id = 3467 then
	sram_write <= x"44446000";
end if;
if first_state_sram_input_id = 3468 then
	sram_write <= x"48622000";
end if;
if first_state_sram_input_id = 3469 then
	sram_write <= x"C89C0000";
end if;
if first_state_sram_input_id = 3470 then
	sram_write <= x"48484000";
end if;
if first_state_sram_input_id = 3471 then
	sram_write <= x"44464000";
end if;
if first_state_sram_input_id = 3472 then
	sram_write <= x"8E04364C";
end if;
if first_state_sram_input_id = 3473 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 3474 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 3475 then
	sram_write <= x"CC3C0028";
end if;
if first_state_sram_input_id = 3476 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 3477 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 3478 then
	sram_write <= x"03DC0038";
end if;
if first_state_sram_input_id = 3479 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 3480 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 3481 then
	sram_write <= x"8200083C";
end if;
if first_state_sram_input_id = 3482 then
	sram_write <= x"07DC0038";
end if;
if first_state_sram_input_id = 3483 then
	sram_write <= x"C03C0018";
end if;
if first_state_sram_input_id = 3484 then
	sram_write <= x"C0220018";
end if;
if first_state_sram_input_id = 3485 then
	sram_write <= x"8220367C";
end if;
if first_state_sram_input_id = 3486 then
	sram_write <= x"82003680";
end if;
if first_state_sram_input_id = 3487 then
	sram_write <= x"44202000";
end if;
if first_state_sram_input_id = 3488 then
	sram_write <= x"022002AC";
end if;
if first_state_sram_input_id = 3489 then
	sram_write <= x"C85C0028";
end if;
if first_state_sram_input_id = 3490 then
	sram_write <= x"44224000";
end if;
if first_state_sram_input_id = 3491 then
	sram_write <= x"C85C0000";
end if;
if first_state_sram_input_id = 3492 then
	sram_write <= x"C43C0030";
end if;
if first_state_sram_input_id = 3493 then
	sram_write <= x"CC3C0038";
end if;
if first_state_sram_input_id = 3494 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 3495 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 3496 then
	sram_write <= x"03DC0048";
end if;
if first_state_sram_input_id = 3497 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 3498 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 3499 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 3500 then
	sram_write <= x"07DC0048";
end if;
if first_state_sram_input_id = 3501 then
	sram_write <= x"C85C0038";
end if;
if first_state_sram_input_id = 3502 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 3503 then
	sram_write <= x"C03C0030";
end if;
if first_state_sram_input_id = 3504 then
	sram_write <= x"CC220000";
end if;
if first_state_sram_input_id = 3505 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 3506 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 3507 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 3508 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 3509 then
	sram_write <= x"028000C8";
end if;
if first_state_sram_input_id = 3510 then
	sram_write <= x"22220220";
end if;
if first_state_sram_input_id = 3511 then
	sram_write <= x"D0282000";
end if;
if first_state_sram_input_id = 3512 then
	sram_write <= x"C8260000";
end if;
if first_state_sram_input_id = 3513 then
	sram_write <= x"C0820014";
end if;
if first_state_sram_input_id = 3514 then
	sram_write <= x"C8480000";
end if;
if first_state_sram_input_id = 3515 then
	sram_write <= x"44224000";
end if;
if first_state_sram_input_id = 3516 then
	sram_write <= x"C8460004";
end if;
if first_state_sram_input_id = 3517 then
	sram_write <= x"C0820014";
end if;
if first_state_sram_input_id = 3518 then
	sram_write <= x"C8680004";
end if;
if first_state_sram_input_id = 3519 then
	sram_write <= x"44446000";
end if;
if first_state_sram_input_id = 3520 then
	sram_write <= x"C8660008";
end if;
if first_state_sram_input_id = 3521 then
	sram_write <= x"C0620014";
end if;
if first_state_sram_input_id = 3522 then
	sram_write <= x"C8860008";
end if;
if first_state_sram_input_id = 3523 then
	sram_write <= x"44668000";
end if;
if first_state_sram_input_id = 3524 then
	sram_write <= x"C0620004";
end if;
if first_state_sram_input_id = 3525 then
	sram_write <= x"02800001";
end if;
if first_state_sram_input_id = 3526 then
	sram_write <= x"826837C8";
end if;
if first_state_sram_input_id = 3527 then
	sram_write <= x"02800002";
end if;
if first_state_sram_input_id = 3528 then
	sram_write <= x"82683728";
end if;
if first_state_sram_input_id = 3529 then
	sram_write <= x"820034A0";
end if;
if first_state_sram_input_id = 3530 then
	sram_write <= x"C0220010";
end if;
if first_state_sram_input_id = 3531 then
	sram_write <= x"C8840000";
end if;
if first_state_sram_input_id = 3532 then
	sram_write <= x"C8A20000";
end if;
if first_state_sram_input_id = 3533 then
	sram_write <= x"4888A000";
end if;
if first_state_sram_input_id = 3534 then
	sram_write <= x"C8A40004";
end if;
if first_state_sram_input_id = 3535 then
	sram_write <= x"C8C20004";
end if;
if first_state_sram_input_id = 3536 then
	sram_write <= x"48AAC000";
end if;
if first_state_sram_input_id = 3537 then
	sram_write <= x"4088A000";
end if;
if first_state_sram_input_id = 3538 then
	sram_write <= x"C8A40008";
end if;
if first_state_sram_input_id = 3539 then
	sram_write <= x"C8C20008";
end if;
if first_state_sram_input_id = 3540 then
	sram_write <= x"48AAC000";
end if;
if first_state_sram_input_id = 3541 then
	sram_write <= x"4088A000";
end if;
if first_state_sram_input_id = 3542 then
	sram_write <= x"8E083764";
end if;
if first_state_sram_input_id = 3543 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 3544 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 3545 then
	sram_write <= x"024002AC";
end if;
if first_state_sram_input_id = 3546 then
	sram_write <= x"C8A20000";
end if;
if first_state_sram_input_id = 3547 then
	sram_write <= x"482A2000";
end if;
if first_state_sram_input_id = 3548 then
	sram_write <= x"C8A20004";
end if;
if first_state_sram_input_id = 3549 then
	sram_write <= x"484A4000";
end if;
if first_state_sram_input_id = 3550 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 3551 then
	sram_write <= x"C8420008";
end if;
if first_state_sram_input_id = 3552 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 3553 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 3554 then
	sram_write <= x"44202000";
end if;
if first_state_sram_input_id = 3555 then
	sram_write <= x"C45C0000";
end if;
if first_state_sram_input_id = 3556 then
	sram_write <= x"CC3C0008";
end if;
if first_state_sram_input_id = 3557 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 3558 then
	sram_write <= x"40208000";
end if;
if first_state_sram_input_id = 3559 then
	sram_write <= x"03DC0018";
end if;
if first_state_sram_input_id = 3560 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 3561 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 3562 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 3563 then
	sram_write <= x"07DC0018";
end if;
if first_state_sram_input_id = 3564 then
	sram_write <= x"C85C0008";
end if;
if first_state_sram_input_id = 3565 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 3566 then
	sram_write <= x"C03C0000";
end if;
if first_state_sram_input_id = 3567 then
	sram_write <= x"CC220000";
end if;
if first_state_sram_input_id = 3568 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 3569 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 3570 then
	sram_write <= x"02600000";
end if;
if first_state_sram_input_id = 3571 then
	sram_write <= x"02800001";
end if;
if first_state_sram_input_id = 3572 then
	sram_write <= x"02A00002";
end if;
if first_state_sram_input_id = 3573 then
	sram_write <= x"CC3C0010";
end if;
if first_state_sram_input_id = 3574 then
	sram_write <= x"CC7C0018";
end if;
if first_state_sram_input_id = 3575 then
	sram_write <= x"CC5C0020";
end if;
if first_state_sram_input_id = 3576 then
	sram_write <= x"C45C0028";
end if;
if first_state_sram_input_id = 3577 then
	sram_write <= x"C43C002C";
end if;
if first_state_sram_input_id = 3578 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 3579 then
	sram_write <= x"03DC0038";
end if;
if first_state_sram_input_id = 3580 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 3581 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 3582 then
	sram_write <= x"8200317C";
end if;
if first_state_sram_input_id = 3583 then
	sram_write <= x"07DC0038";
end if;
if first_state_sram_input_id = 3584 then
	sram_write <= x"8220380C";
end if;
if first_state_sram_input_id = 3585 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 3586 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 3587 then
	sram_write <= x"02600001";
end if;
if first_state_sram_input_id = 3588 then
	sram_write <= x"02800002";
end if;
if first_state_sram_input_id = 3589 then
	sram_write <= x"02A00000";
end if;
if first_state_sram_input_id = 3590 then
	sram_write <= x"C83C0020";
end if;
if first_state_sram_input_id = 3591 then
	sram_write <= x"C85C0018";
end if;
if first_state_sram_input_id = 3592 then
	sram_write <= x"C87C0010";
end if;
if first_state_sram_input_id = 3593 then
	sram_write <= x"C03C002C";
end if;
if first_state_sram_input_id = 3594 then
	sram_write <= x"C05C0028";
end if;
if first_state_sram_input_id = 3595 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 3596 then
	sram_write <= x"03DC0038";
end if;
if first_state_sram_input_id = 3597 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 3598 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 3599 then
	sram_write <= x"8200317C";
end if;
if first_state_sram_input_id = 3600 then
	sram_write <= x"07DC0038";
end if;
if first_state_sram_input_id = 3601 then
	sram_write <= x"82203850";
end if;
if first_state_sram_input_id = 3602 then
	sram_write <= x"02200002";
end if;
if first_state_sram_input_id = 3603 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 3604 then
	sram_write <= x"02600002";
end if;
if first_state_sram_input_id = 3605 then
	sram_write <= x"02800000";
end if;
if first_state_sram_input_id = 3606 then
	sram_write <= x"02A00001";
end if;
if first_state_sram_input_id = 3607 then
	sram_write <= x"C83C0018";
end if;
if first_state_sram_input_id = 3608 then
	sram_write <= x"C85C0010";
end if;
if first_state_sram_input_id = 3609 then
	sram_write <= x"C87C0020";
end if;
if first_state_sram_input_id = 3610 then
	sram_write <= x"C03C002C";
end if;
if first_state_sram_input_id = 3611 then
	sram_write <= x"C05C0028";
end if;
if first_state_sram_input_id = 3612 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 3613 then
	sram_write <= x"03DC0038";
end if;
if first_state_sram_input_id = 3614 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 3615 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 3616 then
	sram_write <= x"8200317C";
end if;
if first_state_sram_input_id = 3617 then
	sram_write <= x"07DC0038";
end if;
if first_state_sram_input_id = 3618 then
	sram_write <= x"82203894";
end if;
if first_state_sram_input_id = 3619 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 3620 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 3621 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 3622 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 3623 then
	sram_write <= x"C8860000";
end if;
if first_state_sram_input_id = 3624 then
	sram_write <= x"44882000";
end if;
if first_state_sram_input_id = 3625 then
	sram_write <= x"C8A60004";
end if;
if first_state_sram_input_id = 3626 then
	sram_write <= x"4888A000";
end if;
if first_state_sram_input_id = 3627 then
	sram_write <= x"C8A40004";
end if;
if first_state_sram_input_id = 3628 then
	sram_write <= x"48A8A000";
end if;
if first_state_sram_input_id = 3629 then
	sram_write <= x"40AA4000";
end if;
if first_state_sram_input_id = 3630 then
	sram_write <= x"8EA038C0";
end if;
if first_state_sram_input_id = 3631 then
	sram_write <= x"820038C4";
end if;
if first_state_sram_input_id = 3632 then
	sram_write <= x"44A0A000";
end if;
if first_state_sram_input_id = 3633 then
	sram_write <= x"C0820010";
end if;
if first_state_sram_input_id = 3634 then
	sram_write <= x"C8C80004";
end if;
if first_state_sram_input_id = 3635 then
	sram_write <= x"8EAC38D8";
end if;
if first_state_sram_input_id = 3636 then
	sram_write <= x"02800000";
end if;
if first_state_sram_input_id = 3637 then
	sram_write <= x"82003918";
end if;
if first_state_sram_input_id = 3638 then
	sram_write <= x"C8A40008";
end if;
if first_state_sram_input_id = 3639 then
	sram_write <= x"48A8A000";
end if;
if first_state_sram_input_id = 3640 then
	sram_write <= x"40AA6000";
end if;
if first_state_sram_input_id = 3641 then
	sram_write <= x"8EA038EC";
end if;
if first_state_sram_input_id = 3642 then
	sram_write <= x"820038F0";
end if;
if first_state_sram_input_id = 3643 then
	sram_write <= x"44A0A000";
end if;
if first_state_sram_input_id = 3644 then
	sram_write <= x"C0820010";
end if;
if first_state_sram_input_id = 3645 then
	sram_write <= x"C8C80008";
end if;
if first_state_sram_input_id = 3646 then
	sram_write <= x"8EAC3904";
end if;
if first_state_sram_input_id = 3647 then
	sram_write <= x"02800000";
end if;
if first_state_sram_input_id = 3648 then
	sram_write <= x"82003918";
end if;
if first_state_sram_input_id = 3649 then
	sram_write <= x"C8A60004";
end if;
if first_state_sram_input_id = 3650 then
	sram_write <= x"8AA03914";
end if;
if first_state_sram_input_id = 3651 then
	sram_write <= x"02800001";
end if;
if first_state_sram_input_id = 3652 then
	sram_write <= x"82003918";
end if;
if first_state_sram_input_id = 3653 then
	sram_write <= x"02800000";
end if;
if first_state_sram_input_id = 3654 then
	sram_write <= x"8280392C";
end if;
if first_state_sram_input_id = 3655 then
	sram_write <= x"022002AC";
end if;
if first_state_sram_input_id = 3656 then
	sram_write <= x"CC820000";
end if;
if first_state_sram_input_id = 3657 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 3658 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 3659 then
	sram_write <= x"C8860008";
end if;
if first_state_sram_input_id = 3660 then
	sram_write <= x"44884000";
end if;
if first_state_sram_input_id = 3661 then
	sram_write <= x"C8A6000C";
end if;
if first_state_sram_input_id = 3662 then
	sram_write <= x"4888A000";
end if;
if first_state_sram_input_id = 3663 then
	sram_write <= x"C8A40000";
end if;
if first_state_sram_input_id = 3664 then
	sram_write <= x"48A8A000";
end if;
if first_state_sram_input_id = 3665 then
	sram_write <= x"40AA2000";
end if;
if first_state_sram_input_id = 3666 then
	sram_write <= x"8EA03950";
end if;
if first_state_sram_input_id = 3667 then
	sram_write <= x"82003954";
end if;
if first_state_sram_input_id = 3668 then
	sram_write <= x"44A0A000";
end if;
if first_state_sram_input_id = 3669 then
	sram_write <= x"C0820010";
end if;
if first_state_sram_input_id = 3670 then
	sram_write <= x"C8C80000";
end if;
if first_state_sram_input_id = 3671 then
	sram_write <= x"8EAC3968";
end if;
if first_state_sram_input_id = 3672 then
	sram_write <= x"02800000";
end if;
if first_state_sram_input_id = 3673 then
	sram_write <= x"820039A8";
end if;
if first_state_sram_input_id = 3674 then
	sram_write <= x"C8A40008";
end if;
if first_state_sram_input_id = 3675 then
	sram_write <= x"48A8A000";
end if;
if first_state_sram_input_id = 3676 then
	sram_write <= x"40AA6000";
end if;
if first_state_sram_input_id = 3677 then
	sram_write <= x"8EA0397C";
end if;
if first_state_sram_input_id = 3678 then
	sram_write <= x"82003980";
end if;
if first_state_sram_input_id = 3679 then
	sram_write <= x"44A0A000";
end if;
if first_state_sram_input_id = 3680 then
	sram_write <= x"C0820010";
end if;
if first_state_sram_input_id = 3681 then
	sram_write <= x"C8C80008";
end if;
if first_state_sram_input_id = 3682 then
	sram_write <= x"8EAC3994";
end if;
if first_state_sram_input_id = 3683 then
	sram_write <= x"02800000";
end if;
if first_state_sram_input_id = 3684 then
	sram_write <= x"820039A8";
end if;
if first_state_sram_input_id = 3685 then
	sram_write <= x"C8A6000C";
end if;
if first_state_sram_input_id = 3686 then
	sram_write <= x"8AA039A4";
end if;
if first_state_sram_input_id = 3687 then
	sram_write <= x"02800001";
end if;
if first_state_sram_input_id = 3688 then
	sram_write <= x"820039A8";
end if;
if first_state_sram_input_id = 3689 then
	sram_write <= x"02800000";
end if;
if first_state_sram_input_id = 3690 then
	sram_write <= x"828039BC";
end if;
if first_state_sram_input_id = 3691 then
	sram_write <= x"022002AC";
end if;
if first_state_sram_input_id = 3692 then
	sram_write <= x"CC820000";
end if;
if first_state_sram_input_id = 3693 then
	sram_write <= x"02200002";
end if;
if first_state_sram_input_id = 3694 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 3695 then
	sram_write <= x"C8860010";
end if;
if first_state_sram_input_id = 3696 then
	sram_write <= x"44686000";
end if;
if first_state_sram_input_id = 3697 then
	sram_write <= x"C8860014";
end if;
if first_state_sram_input_id = 3698 then
	sram_write <= x"48668000";
end if;
if first_state_sram_input_id = 3699 then
	sram_write <= x"C8840000";
end if;
if first_state_sram_input_id = 3700 then
	sram_write <= x"48868000";
end if;
if first_state_sram_input_id = 3701 then
	sram_write <= x"40282000";
end if;
if first_state_sram_input_id = 3702 then
	sram_write <= x"8E2039E0";
end if;
if first_state_sram_input_id = 3703 then
	sram_write <= x"820039E4";
end if;
if first_state_sram_input_id = 3704 then
	sram_write <= x"44202000";
end if;
if first_state_sram_input_id = 3705 then
	sram_write <= x"C0820010";
end if;
if first_state_sram_input_id = 3706 then
	sram_write <= x"C8880000";
end if;
if first_state_sram_input_id = 3707 then
	sram_write <= x"8E2839F8";
end if;
if first_state_sram_input_id = 3708 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 3709 then
	sram_write <= x"82003A38";
end if;
if first_state_sram_input_id = 3710 then
	sram_write <= x"C8240004";
end if;
if first_state_sram_input_id = 3711 then
	sram_write <= x"48262000";
end if;
if first_state_sram_input_id = 3712 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 3713 then
	sram_write <= x"8E203A0C";
end if;
if first_state_sram_input_id = 3714 then
	sram_write <= x"82003A10";
end if;
if first_state_sram_input_id = 3715 then
	sram_write <= x"44202000";
end if;
if first_state_sram_input_id = 3716 then
	sram_write <= x"C0220010";
end if;
if first_state_sram_input_id = 3717 then
	sram_write <= x"C8420004";
end if;
if first_state_sram_input_id = 3718 then
	sram_write <= x"8E243A24";
end if;
if first_state_sram_input_id = 3719 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 3720 then
	sram_write <= x"82003A38";
end if;
if first_state_sram_input_id = 3721 then
	sram_write <= x"C8260014";
end if;
if first_state_sram_input_id = 3722 then
	sram_write <= x"8A203A34";
end if;
if first_state_sram_input_id = 3723 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 3724 then
	sram_write <= x"82003A38";
end if;
if first_state_sram_input_id = 3725 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 3726 then
	sram_write <= x"82203A4C";
end if;
if first_state_sram_input_id = 3727 then
	sram_write <= x"022002AC";
end if;
if first_state_sram_input_id = 3728 then
	sram_write <= x"CC620000";
end if;
if first_state_sram_input_id = 3729 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 3730 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 3731 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 3732 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 3733 then
	sram_write <= x"C8840000";
end if;
if first_state_sram_input_id = 3734 then
	sram_write <= x"8A803BCC";
end if;
if first_state_sram_input_id = 3735 then
	sram_write <= x"C8A40004";
end if;
if first_state_sram_input_id = 3736 then
	sram_write <= x"48AA2000";
end if;
if first_state_sram_input_id = 3737 then
	sram_write <= x"C8C40008";
end if;
if first_state_sram_input_id = 3738 then
	sram_write <= x"48CC4000";
end if;
if first_state_sram_input_id = 3739 then
	sram_write <= x"40AAC000";
end if;
if first_state_sram_input_id = 3740 then
	sram_write <= x"C8C4000C";
end if;
if first_state_sram_input_id = 3741 then
	sram_write <= x"48CC6000";
end if;
if first_state_sram_input_id = 3742 then
	sram_write <= x"40AAC000";
end if;
if first_state_sram_input_id = 3743 then
	sram_write <= x"48C22000";
end if;
if first_state_sram_input_id = 3744 then
	sram_write <= x"C0620010";
end if;
if first_state_sram_input_id = 3745 then
	sram_write <= x"C8E60000";
end if;
if first_state_sram_input_id = 3746 then
	sram_write <= x"48CCE000";
end if;
if first_state_sram_input_id = 3747 then
	sram_write <= x"48E44000";
end if;
if first_state_sram_input_id = 3748 then
	sram_write <= x"C0620010";
end if;
if first_state_sram_input_id = 3749 then
	sram_write <= x"C9060004";
end if;
if first_state_sram_input_id = 3750 then
	sram_write <= x"48EF0000";
end if;
if first_state_sram_input_id = 3751 then
	sram_write <= x"40CCE000";
end if;
if first_state_sram_input_id = 3752 then
	sram_write <= x"48E66000";
end if;
if first_state_sram_input_id = 3753 then
	sram_write <= x"C0620010";
end if;
if first_state_sram_input_id = 3754 then
	sram_write <= x"C9060008";
end if;
if first_state_sram_input_id = 3755 then
	sram_write <= x"48EF0000";
end if;
if first_state_sram_input_id = 3756 then
	sram_write <= x"40CCE000";
end if;
if first_state_sram_input_id = 3757 then
	sram_write <= x"C062000C";
end if;
if first_state_sram_input_id = 3758 then
	sram_write <= x"82603AFC";
end if;
if first_state_sram_input_id = 3759 then
	sram_write <= x"48E46000";
end if;
if first_state_sram_input_id = 3760 then
	sram_write <= x"C0620024";
end if;
if first_state_sram_input_id = 3761 then
	sram_write <= x"C9060000";
end if;
if first_state_sram_input_id = 3762 then
	sram_write <= x"48EF0000";
end if;
if first_state_sram_input_id = 3763 then
	sram_write <= x"40CCE000";
end if;
if first_state_sram_input_id = 3764 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 3765 then
	sram_write <= x"C0620024";
end if;
if first_state_sram_input_id = 3766 then
	sram_write <= x"C8E60004";
end if;
if first_state_sram_input_id = 3767 then
	sram_write <= x"4866E000";
end if;
if first_state_sram_input_id = 3768 then
	sram_write <= x"406C6000";
end if;
if first_state_sram_input_id = 3769 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 3770 then
	sram_write <= x"C0620024";
end if;
if first_state_sram_input_id = 3771 then
	sram_write <= x"C8460008";
end if;
if first_state_sram_input_id = 3772 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 3773 then
	sram_write <= x"40262000";
end if;
if first_state_sram_input_id = 3774 then
	sram_write <= x"82003B00";
end if;
if first_state_sram_input_id = 3775 then
	sram_write <= x"4020C000";
end if;
if first_state_sram_input_id = 3776 then
	sram_write <= x"C0620004";
end if;
if first_state_sram_input_id = 3777 then
	sram_write <= x"02800003";
end if;
if first_state_sram_input_id = 3778 then
	sram_write <= x"82683B10";
end if;
if first_state_sram_input_id = 3779 then
	sram_write <= x"82003B18";
end if;
if first_state_sram_input_id = 3780 then
	sram_write <= x"C84000A8";
end if;
if first_state_sram_input_id = 3781 then
	sram_write <= x"44224000";
end if;
if first_state_sram_input_id = 3782 then
	sram_write <= x"484AA000";
end if;
if first_state_sram_input_id = 3783 then
	sram_write <= x"48282000";
end if;
if first_state_sram_input_id = 3784 then
	sram_write <= x"44242000";
end if;
if first_state_sram_input_id = 3785 then
	sram_write <= x"8E023B30";
end if;
if first_state_sram_input_id = 3786 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 3787 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 3788 then
	sram_write <= x"C0220018";
end if;
if first_state_sram_input_id = 3789 then
	sram_write <= x"82203B80";
end if;
if first_state_sram_input_id = 3790 then
	sram_write <= x"022002AC";
end if;
if first_state_sram_input_id = 3791 then
	sram_write <= x"C43C0000";
end if;
if first_state_sram_input_id = 3792 then
	sram_write <= x"C45C0004";
end if;
if first_state_sram_input_id = 3793 then
	sram_write <= x"CCBC0008";
end if;
if first_state_sram_input_id = 3794 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 3795 then
	sram_write <= x"03DC0018";
end if;
if first_state_sram_input_id = 3796 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 3797 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 3798 then
	sram_write <= x"8200083C";
end if;
if first_state_sram_input_id = 3799 then
	sram_write <= x"07DC0018";
end if;
if first_state_sram_input_id = 3800 then
	sram_write <= x"C85C0008";
end if;
if first_state_sram_input_id = 3801 then
	sram_write <= x"40242000";
end if;
if first_state_sram_input_id = 3802 then
	sram_write <= x"C03C0004";
end if;
if first_state_sram_input_id = 3803 then
	sram_write <= x"C8420010";
end if;
if first_state_sram_input_id = 3804 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 3805 then
	sram_write <= x"C03C0000";
end if;
if first_state_sram_input_id = 3806 then
	sram_write <= x"CC220000";
end if;
if first_state_sram_input_id = 3807 then
	sram_write <= x"82003BC4";
end if;
if first_state_sram_input_id = 3808 then
	sram_write <= x"022002AC";
end if;
if first_state_sram_input_id = 3809 then
	sram_write <= x"C43C0010";
end if;
if first_state_sram_input_id = 3810 then
	sram_write <= x"C45C0004";
end if;
if first_state_sram_input_id = 3811 then
	sram_write <= x"CCBC0008";
end if;
if first_state_sram_input_id = 3812 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 3813 then
	sram_write <= x"03DC001C";
end if;
if first_state_sram_input_id = 3814 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 3815 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 3816 then
	sram_write <= x"8200083C";
end if;
if first_state_sram_input_id = 3817 then
	sram_write <= x"07DC001C";
end if;
if first_state_sram_input_id = 3818 then
	sram_write <= x"C85C0008";
end if;
if first_state_sram_input_id = 3819 then
	sram_write <= x"44242000";
end if;
if first_state_sram_input_id = 3820 then
	sram_write <= x"C03C0004";
end if;
if first_state_sram_input_id = 3821 then
	sram_write <= x"C8420010";
end if;
if first_state_sram_input_id = 3822 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 3823 then
	sram_write <= x"C03C0010";
end if;
if first_state_sram_input_id = 3824 then
	sram_write <= x"CC220000";
end if;
if first_state_sram_input_id = 3825 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 3826 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 3827 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 3828 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 3829 then
	sram_write <= x"C8840000";
end if;
if first_state_sram_input_id = 3830 then
	sram_write <= x"8A803CBC";
end if;
if first_state_sram_input_id = 3831 then
	sram_write <= x"C8A40004";
end if;
if first_state_sram_input_id = 3832 then
	sram_write <= x"482A2000";
end if;
if first_state_sram_input_id = 3833 then
	sram_write <= x"C8A40008";
end if;
if first_state_sram_input_id = 3834 then
	sram_write <= x"484A4000";
end if;
if first_state_sram_input_id = 3835 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 3836 then
	sram_write <= x"C844000C";
end if;
if first_state_sram_input_id = 3837 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 3838 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 3839 then
	sram_write <= x"C846000C";
end if;
if first_state_sram_input_id = 3840 then
	sram_write <= x"48622000";
end if;
if first_state_sram_input_id = 3841 then
	sram_write <= x"48484000";
end if;
if first_state_sram_input_id = 3842 then
	sram_write <= x"44464000";
end if;
if first_state_sram_input_id = 3843 then
	sram_write <= x"8E043C18";
end if;
if first_state_sram_input_id = 3844 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 3845 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 3846 then
	sram_write <= x"C0220018";
end if;
if first_state_sram_input_id = 3847 then
	sram_write <= x"82203C6C";
end if;
if first_state_sram_input_id = 3848 then
	sram_write <= x"022002AC";
end if;
if first_state_sram_input_id = 3849 then
	sram_write <= x"C43C0000";
end if;
if first_state_sram_input_id = 3850 then
	sram_write <= x"C45C0004";
end if;
if first_state_sram_input_id = 3851 then
	sram_write <= x"CC3C0008";
end if;
if first_state_sram_input_id = 3852 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 3853 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 3854 then
	sram_write <= x"03DC0018";
end if;
if first_state_sram_input_id = 3855 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 3856 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 3857 then
	sram_write <= x"8200083C";
end if;
if first_state_sram_input_id = 3858 then
	sram_write <= x"07DC0018";
end if;
if first_state_sram_input_id = 3859 then
	sram_write <= x"C85C0008";
end if;
if first_state_sram_input_id = 3860 then
	sram_write <= x"40242000";
end if;
if first_state_sram_input_id = 3861 then
	sram_write <= x"C03C0004";
end if;
if first_state_sram_input_id = 3862 then
	sram_write <= x"C8420010";
end if;
if first_state_sram_input_id = 3863 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 3864 then
	sram_write <= x"C03C0000";
end if;
if first_state_sram_input_id = 3865 then
	sram_write <= x"CC220000";
end if;
if first_state_sram_input_id = 3866 then
	sram_write <= x"82003CB4";
end if;
if first_state_sram_input_id = 3867 then
	sram_write <= x"022002AC";
end if;
if first_state_sram_input_id = 3868 then
	sram_write <= x"C43C0010";
end if;
if first_state_sram_input_id = 3869 then
	sram_write <= x"C45C0004";
end if;
if first_state_sram_input_id = 3870 then
	sram_write <= x"CC3C0008";
end if;
if first_state_sram_input_id = 3871 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 3872 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 3873 then
	sram_write <= x"03DC001C";
end if;
if first_state_sram_input_id = 3874 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 3875 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 3876 then
	sram_write <= x"8200083C";
end if;
if first_state_sram_input_id = 3877 then
	sram_write <= x"07DC001C";
end if;
if first_state_sram_input_id = 3878 then
	sram_write <= x"C85C0008";
end if;
if first_state_sram_input_id = 3879 then
	sram_write <= x"44242000";
end if;
if first_state_sram_input_id = 3880 then
	sram_write <= x"C03C0004";
end if;
if first_state_sram_input_id = 3881 then
	sram_write <= x"C8420010";
end if;
if first_state_sram_input_id = 3882 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 3883 then
	sram_write <= x"C03C0010";
end if;
if first_state_sram_input_id = 3884 then
	sram_write <= x"CC220000";
end if;
if first_state_sram_input_id = 3885 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 3886 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 3887 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 3888 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 3889 then
	sram_write <= x"02600006";
end if;
if first_state_sram_input_id = 3890 then
	sram_write <= x"40200000";
end if;
if first_state_sram_input_id = 3891 then
	sram_write <= x"C45C0000";
end if;
if first_state_sram_input_id = 3892 then
	sram_write <= x"C43C0004";
end if;
if first_state_sram_input_id = 3893 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 3894 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 3895 then
	sram_write <= x"03DC0010";
end if;
if first_state_sram_input_id = 3896 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 3897 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 3898 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 3899 then
	sram_write <= x"07DC0010";
end if;
if first_state_sram_input_id = 3900 then
	sram_write <= x"C05C0004";
end if;
if first_state_sram_input_id = 3901 then
	sram_write <= x"C8240000";
end if;
if first_state_sram_input_id = 3902 then
	sram_write <= x"8A203D78";
end if;
if first_state_sram_input_id = 3903 then
	sram_write <= x"C07C0000";
end if;
if first_state_sram_input_id = 3904 then
	sram_write <= x"C0860018";
end if;
if first_state_sram_input_id = 3905 then
	sram_write <= x"C8240000";
end if;
if first_state_sram_input_id = 3906 then
	sram_write <= x"8E203D14";
end if;
if first_state_sram_input_id = 3907 then
	sram_write <= x"02A00000";
end if;
if first_state_sram_input_id = 3908 then
	sram_write <= x"82003D18";
end if;
if first_state_sram_input_id = 3909 then
	sram_write <= x"02A00001";
end if;
if first_state_sram_input_id = 3910 then
	sram_write <= x"82803D30";
end if;
if first_state_sram_input_id = 3911 then
	sram_write <= x"8E203D28";
end if;
if first_state_sram_input_id = 3912 then
	sram_write <= x"02800001";
end if;
if first_state_sram_input_id = 3913 then
	sram_write <= x"82003D2C";
end if;
if first_state_sram_input_id = 3914 then
	sram_write <= x"02800000";
end if;
if first_state_sram_input_id = 3915 then
	sram_write <= x"82003D34";
end if;
if first_state_sram_input_id = 3916 then
	sram_write <= x"008A0000";
end if;
if first_state_sram_input_id = 3917 then
	sram_write <= x"C0A60010";
end if;
if first_state_sram_input_id = 3918 then
	sram_write <= x"C82A0000";
end if;
if first_state_sram_input_id = 3919 then
	sram_write <= x"82803D44";
end if;
if first_state_sram_input_id = 3920 then
	sram_write <= x"82003D48";
end if;
if first_state_sram_input_id = 3921 then
	sram_write <= x"44202000";
end if;
if first_state_sram_input_id = 3922 then
	sram_write <= x"CC220000";
end if;
if first_state_sram_input_id = 3923 then
	sram_write <= x"C8240000";
end if;
if first_state_sram_input_id = 3924 then
	sram_write <= x"C43C0008";
end if;
if first_state_sram_input_id = 3925 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 3926 then
	sram_write <= x"03DC0014";
end if;
if first_state_sram_input_id = 3927 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 3928 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 3929 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 3930 then
	sram_write <= x"07DC0014";
end if;
if first_state_sram_input_id = 3931 then
	sram_write <= x"C03C0008";
end if;
if first_state_sram_input_id = 3932 then
	sram_write <= x"CC220004";
end if;
if first_state_sram_input_id = 3933 then
	sram_write <= x"82003D7C";
end if;
if first_state_sram_input_id = 3934 then
	sram_write <= x"CC020004";
end if;
if first_state_sram_input_id = 3935 then
	sram_write <= x"C05C0004";
end if;
if first_state_sram_input_id = 3936 then
	sram_write <= x"C8240004";
end if;
if first_state_sram_input_id = 3937 then
	sram_write <= x"8A203E04";
end if;
if first_state_sram_input_id = 3938 then
	sram_write <= x"C07C0000";
end if;
if first_state_sram_input_id = 3939 then
	sram_write <= x"C0860018";
end if;
if first_state_sram_input_id = 3940 then
	sram_write <= x"C8240004";
end if;
if first_state_sram_input_id = 3941 then
	sram_write <= x"8E203DA0";
end if;
if first_state_sram_input_id = 3942 then
	sram_write <= x"02A00000";
end if;
if first_state_sram_input_id = 3943 then
	sram_write <= x"82003DA4";
end if;
if first_state_sram_input_id = 3944 then
	sram_write <= x"02A00001";
end if;
if first_state_sram_input_id = 3945 then
	sram_write <= x"82803DBC";
end if;
if first_state_sram_input_id = 3946 then
	sram_write <= x"8E203DB4";
end if;
if first_state_sram_input_id = 3947 then
	sram_write <= x"02800001";
end if;
if first_state_sram_input_id = 3948 then
	sram_write <= x"82003DB8";
end if;
if first_state_sram_input_id = 3949 then
	sram_write <= x"02800000";
end if;
if first_state_sram_input_id = 3950 then
	sram_write <= x"82003DC0";
end if;
if first_state_sram_input_id = 3951 then
	sram_write <= x"008A0000";
end if;
if first_state_sram_input_id = 3952 then
	sram_write <= x"C0A60010";
end if;
if first_state_sram_input_id = 3953 then
	sram_write <= x"C82A0004";
end if;
if first_state_sram_input_id = 3954 then
	sram_write <= x"82803DD0";
end if;
if first_state_sram_input_id = 3955 then
	sram_write <= x"82003DD4";
end if;
if first_state_sram_input_id = 3956 then
	sram_write <= x"44202000";
end if;
if first_state_sram_input_id = 3957 then
	sram_write <= x"CC220008";
end if;
if first_state_sram_input_id = 3958 then
	sram_write <= x"C8240004";
end if;
if first_state_sram_input_id = 3959 then
	sram_write <= x"C43C0008";
end if;
if first_state_sram_input_id = 3960 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 3961 then
	sram_write <= x"03DC0014";
end if;
if first_state_sram_input_id = 3962 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 3963 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 3964 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 3965 then
	sram_write <= x"07DC0014";
end if;
if first_state_sram_input_id = 3966 then
	sram_write <= x"C03C0008";
end if;
if first_state_sram_input_id = 3967 then
	sram_write <= x"CC22000C";
end if;
if first_state_sram_input_id = 3968 then
	sram_write <= x"82003E08";
end if;
if first_state_sram_input_id = 3969 then
	sram_write <= x"CC02000C";
end if;
if first_state_sram_input_id = 3970 then
	sram_write <= x"C05C0004";
end if;
if first_state_sram_input_id = 3971 then
	sram_write <= x"C8240008";
end if;
if first_state_sram_input_id = 3972 then
	sram_write <= x"8A203E90";
end if;
if first_state_sram_input_id = 3973 then
	sram_write <= x"C07C0000";
end if;
if first_state_sram_input_id = 3974 then
	sram_write <= x"C0860018";
end if;
if first_state_sram_input_id = 3975 then
	sram_write <= x"C8240008";
end if;
if first_state_sram_input_id = 3976 then
	sram_write <= x"8E203E2C";
end if;
if first_state_sram_input_id = 3977 then
	sram_write <= x"02A00000";
end if;
if first_state_sram_input_id = 3978 then
	sram_write <= x"82003E30";
end if;
if first_state_sram_input_id = 3979 then
	sram_write <= x"02A00001";
end if;
if first_state_sram_input_id = 3980 then
	sram_write <= x"82803E48";
end if;
if first_state_sram_input_id = 3981 then
	sram_write <= x"8E203E40";
end if;
if first_state_sram_input_id = 3982 then
	sram_write <= x"02800001";
end if;
if first_state_sram_input_id = 3983 then
	sram_write <= x"82003E44";
end if;
if first_state_sram_input_id = 3984 then
	sram_write <= x"02800000";
end if;
if first_state_sram_input_id = 3985 then
	sram_write <= x"82003E4C";
end if;
if first_state_sram_input_id = 3986 then
	sram_write <= x"008A0000";
end if;
if first_state_sram_input_id = 3987 then
	sram_write <= x"C0660010";
end if;
if first_state_sram_input_id = 3988 then
	sram_write <= x"C8260008";
end if;
if first_state_sram_input_id = 3989 then
	sram_write <= x"82803E5C";
end if;
if first_state_sram_input_id = 3990 then
	sram_write <= x"82003E60";
end if;
if first_state_sram_input_id = 3991 then
	sram_write <= x"44202000";
end if;
if first_state_sram_input_id = 3992 then
	sram_write <= x"CC220010";
end if;
if first_state_sram_input_id = 3993 then
	sram_write <= x"C8240008";
end if;
if first_state_sram_input_id = 3994 then
	sram_write <= x"C43C0008";
end if;
if first_state_sram_input_id = 3995 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 3996 then
	sram_write <= x"03DC0014";
end if;
if first_state_sram_input_id = 3997 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 3998 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 3999 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 4000 then
	sram_write <= x"07DC0014";
end if;
if first_state_sram_input_id = 4001 then
	sram_write <= x"C03C0008";
end if;
if first_state_sram_input_id = 4002 then
	sram_write <= x"CC220014";
end if;
if first_state_sram_input_id = 4003 then
	sram_write <= x"82003E94";
end if;
if first_state_sram_input_id = 4004 then
	sram_write <= x"CC020014";
end if;
if first_state_sram_input_id = 4005 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 4006 then
	sram_write <= x"02600004";
end if;
if first_state_sram_input_id = 4007 then
	sram_write <= x"40200000";
end if;
if first_state_sram_input_id = 4008 then
	sram_write <= x"C45C0000";
end if;
if first_state_sram_input_id = 4009 then
	sram_write <= x"C43C0004";
end if;
if first_state_sram_input_id = 4010 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 4011 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 4012 then
	sram_write <= x"03DC0010";
end if;
if first_state_sram_input_id = 4013 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 4014 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 4015 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 4016 then
	sram_write <= x"07DC0010";
end if;
if first_state_sram_input_id = 4017 then
	sram_write <= x"C05C0004";
end if;
if first_state_sram_input_id = 4018 then
	sram_write <= x"C8240000";
end if;
if first_state_sram_input_id = 4019 then
	sram_write <= x"C07C0000";
end if;
if first_state_sram_input_id = 4020 then
	sram_write <= x"C0860010";
end if;
if first_state_sram_input_id = 4021 then
	sram_write <= x"C8480000";
end if;
if first_state_sram_input_id = 4022 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 4023 then
	sram_write <= x"C8440004";
end if;
if first_state_sram_input_id = 4024 then
	sram_write <= x"C0860010";
end if;
if first_state_sram_input_id = 4025 then
	sram_write <= x"C8680004";
end if;
if first_state_sram_input_id = 4026 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 4027 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 4028 then
	sram_write <= x"C8440008";
end if;
if first_state_sram_input_id = 4029 then
	sram_write <= x"C0460010";
end if;
if first_state_sram_input_id = 4030 then
	sram_write <= x"C8640008";
end if;
if first_state_sram_input_id = 4031 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 4032 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 4033 then
	sram_write <= x"8E023F10";
end if;
if first_state_sram_input_id = 4034 then
	sram_write <= x"CC020000";
end if;
if first_state_sram_input_id = 4035 then
	sram_write <= x"82004008";
end if;
if first_state_sram_input_id = 4036 then
	sram_write <= x"CC3C0008";
end if;
if first_state_sram_input_id = 4037 then
	sram_write <= x"C43C0010";
end if;
if first_state_sram_input_id = 4038 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 4039 then
	sram_write <= x"03DC001C";
end if;
if first_state_sram_input_id = 4040 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 4041 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 4042 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 4043 then
	sram_write <= x"07DC001C";
end if;
if first_state_sram_input_id = 4044 then
	sram_write <= x"44202000";
end if;
if first_state_sram_input_id = 4045 then
	sram_write <= x"C03C0010";
end if;
if first_state_sram_input_id = 4046 then
	sram_write <= x"CC220000";
end if;
if first_state_sram_input_id = 4047 then
	sram_write <= x"C05C0000";
end if;
if first_state_sram_input_id = 4048 then
	sram_write <= x"C0640010";
end if;
if first_state_sram_input_id = 4049 then
	sram_write <= x"C8260000";
end if;
if first_state_sram_input_id = 4050 then
	sram_write <= x"C85C0008";
end if;
if first_state_sram_input_id = 4051 then
	sram_write <= x"CC3C0018";
end if;
if first_state_sram_input_id = 4052 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 4053 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 4054 then
	sram_write <= x"03DC0028";
end if;
if first_state_sram_input_id = 4055 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 4056 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 4057 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 4058 then
	sram_write <= x"07DC0028";
end if;
if first_state_sram_input_id = 4059 then
	sram_write <= x"C85C0018";
end if;
if first_state_sram_input_id = 4060 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 4061 then
	sram_write <= x"44202000";
end if;
if first_state_sram_input_id = 4062 then
	sram_write <= x"C03C0010";
end if;
if first_state_sram_input_id = 4063 then
	sram_write <= x"CC220004";
end if;
if first_state_sram_input_id = 4064 then
	sram_write <= x"C05C0000";
end if;
if first_state_sram_input_id = 4065 then
	sram_write <= x"C0640010";
end if;
if first_state_sram_input_id = 4066 then
	sram_write <= x"C8260004";
end if;
if first_state_sram_input_id = 4067 then
	sram_write <= x"C85C0008";
end if;
if first_state_sram_input_id = 4068 then
	sram_write <= x"CC3C0020";
end if;
if first_state_sram_input_id = 4069 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 4070 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 4071 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 4072 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 4073 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 4074 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 4075 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 4076 then
	sram_write <= x"C85C0020";
end if;
if first_state_sram_input_id = 4077 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 4078 then
	sram_write <= x"44202000";
end if;
if first_state_sram_input_id = 4079 then
	sram_write <= x"C03C0010";
end if;
if first_state_sram_input_id = 4080 then
	sram_write <= x"CC220008";
end if;
if first_state_sram_input_id = 4081 then
	sram_write <= x"C05C0000";
end if;
if first_state_sram_input_id = 4082 then
	sram_write <= x"C0440010";
end if;
if first_state_sram_input_id = 4083 then
	sram_write <= x"C8240008";
end if;
if first_state_sram_input_id = 4084 then
	sram_write <= x"C85C0008";
end if;
if first_state_sram_input_id = 4085 then
	sram_write <= x"CC3C0028";
end if;
if first_state_sram_input_id = 4086 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 4087 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 4088 then
	sram_write <= x"03DC0038";
end if;
if first_state_sram_input_id = 4089 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 4090 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 4091 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 4092 then
	sram_write <= x"07DC0038";
end if;
if first_state_sram_input_id = 4093 then
	sram_write <= x"C85C0028";
end if;
if first_state_sram_input_id = 4094 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 4095 then
	sram_write <= x"44202000";
end if;
if first_state_sram_input_id = 4096 then
	sram_write <= x"C03C0010";
end if;
if first_state_sram_input_id = 4097 then
	sram_write <= x"CC22000C";
end if;
if first_state_sram_input_id = 4098 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 4099 then
	sram_write <= x"02600005";
end if;
if first_state_sram_input_id = 4100 then
	sram_write <= x"40200000";
end if;
if first_state_sram_input_id = 4101 then
	sram_write <= x"C45C0000";
end if;
if first_state_sram_input_id = 4102 then
	sram_write <= x"C43C0004";
end if;
if first_state_sram_input_id = 4103 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 4104 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 4105 then
	sram_write <= x"03DC0010";
end if;
if first_state_sram_input_id = 4106 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 4107 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 4108 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 4109 then
	sram_write <= x"07DC0010";
end if;
if first_state_sram_input_id = 4110 then
	sram_write <= x"C05C0004";
end if;
if first_state_sram_input_id = 4111 then
	sram_write <= x"C8240000";
end if;
if first_state_sram_input_id = 4112 then
	sram_write <= x"C8440004";
end if;
if first_state_sram_input_id = 4113 then
	sram_write <= x"C8640008";
end if;
if first_state_sram_input_id = 4114 then
	sram_write <= x"48822000";
end if;
if first_state_sram_input_id = 4115 then
	sram_write <= x"C07C0000";
end if;
if first_state_sram_input_id = 4116 then
	sram_write <= x"C0860010";
end if;
if first_state_sram_input_id = 4117 then
	sram_write <= x"C8A80000";
end if;
if first_state_sram_input_id = 4118 then
	sram_write <= x"4888A000";
end if;
if first_state_sram_input_id = 4119 then
	sram_write <= x"48A44000";
end if;
if first_state_sram_input_id = 4120 then
	sram_write <= x"C0860010";
end if;
if first_state_sram_input_id = 4121 then
	sram_write <= x"C8C80004";
end if;
if first_state_sram_input_id = 4122 then
	sram_write <= x"48AAC000";
end if;
if first_state_sram_input_id = 4123 then
	sram_write <= x"4088A000";
end if;
if first_state_sram_input_id = 4124 then
	sram_write <= x"48A66000";
end if;
if first_state_sram_input_id = 4125 then
	sram_write <= x"C0860010";
end if;
if first_state_sram_input_id = 4126 then
	sram_write <= x"C8C80008";
end if;
if first_state_sram_input_id = 4127 then
	sram_write <= x"48AAC000";
end if;
if first_state_sram_input_id = 4128 then
	sram_write <= x"4088A000";
end if;
if first_state_sram_input_id = 4129 then
	sram_write <= x"C086000C";
end if;
if first_state_sram_input_id = 4130 then
	sram_write <= x"828040CC";
end if;
if first_state_sram_input_id = 4131 then
	sram_write <= x"48A46000";
end if;
if first_state_sram_input_id = 4132 then
	sram_write <= x"C0860024";
end if;
if first_state_sram_input_id = 4133 then
	sram_write <= x"C8C80000";
end if;
if first_state_sram_input_id = 4134 then
	sram_write <= x"48AAC000";
end if;
if first_state_sram_input_id = 4135 then
	sram_write <= x"4088A000";
end if;
if first_state_sram_input_id = 4136 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 4137 then
	sram_write <= x"C0860024";
end if;
if first_state_sram_input_id = 4138 then
	sram_write <= x"C8A80004";
end if;
if first_state_sram_input_id = 4139 then
	sram_write <= x"4866A000";
end if;
if first_state_sram_input_id = 4140 then
	sram_write <= x"40686000";
end if;
if first_state_sram_input_id = 4141 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 4142 then
	sram_write <= x"C0860024";
end if;
if first_state_sram_input_id = 4143 then
	sram_write <= x"C8480008";
end if;
if first_state_sram_input_id = 4144 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 4145 then
	sram_write <= x"40262000";
end if;
if first_state_sram_input_id = 4146 then
	sram_write <= x"820040D0";
end if;
if first_state_sram_input_id = 4147 then
	sram_write <= x"40208000";
end if;
if first_state_sram_input_id = 4148 then
	sram_write <= x"C8440000";
end if;
if first_state_sram_input_id = 4149 then
	sram_write <= x"C0860010";
end if;
if first_state_sram_input_id = 4150 then
	sram_write <= x"C8680000";
end if;
if first_state_sram_input_id = 4151 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 4152 then
	sram_write <= x"44404000";
end if;
if first_state_sram_input_id = 4153 then
	sram_write <= x"C8640004";
end if;
if first_state_sram_input_id = 4154 then
	sram_write <= x"C0860010";
end if;
if first_state_sram_input_id = 4155 then
	sram_write <= x"C8880004";
end if;
if first_state_sram_input_id = 4156 then
	sram_write <= x"48668000";
end if;
if first_state_sram_input_id = 4157 then
	sram_write <= x"44606000";
end if;
if first_state_sram_input_id = 4158 then
	sram_write <= x"C8840008";
end if;
if first_state_sram_input_id = 4159 then
	sram_write <= x"C0860010";
end if;
if first_state_sram_input_id = 4160 then
	sram_write <= x"C8A80008";
end if;
if first_state_sram_input_id = 4161 then
	sram_write <= x"4888A000";
end if;
if first_state_sram_input_id = 4162 then
	sram_write <= x"44808000";
end if;
if first_state_sram_input_id = 4163 then
	sram_write <= x"CC220000";
end if;
if first_state_sram_input_id = 4164 then
	sram_write <= x"C086000C";
end if;
if first_state_sram_input_id = 4165 then
	sram_write <= x"CC3C0008";
end if;
if first_state_sram_input_id = 4166 then
	sram_write <= x"82804264";
end if;
if first_state_sram_input_id = 4167 then
	sram_write <= x"C8A40008";
end if;
if first_state_sram_input_id = 4168 then
	sram_write <= x"C0860024";
end if;
if first_state_sram_input_id = 4169 then
	sram_write <= x"C8C80004";
end if;
if first_state_sram_input_id = 4170 then
	sram_write <= x"48AAC000";
end if;
if first_state_sram_input_id = 4171 then
	sram_write <= x"C8C40004";
end if;
if first_state_sram_input_id = 4172 then
	sram_write <= x"C0860024";
end if;
if first_state_sram_input_id = 4173 then
	sram_write <= x"C8E80008";
end if;
if first_state_sram_input_id = 4174 then
	sram_write <= x"48CCE000";
end if;
if first_state_sram_input_id = 4175 then
	sram_write <= x"40AAC000";
end if;
if first_state_sram_input_id = 4176 then
	sram_write <= x"C8C00080";
end if;
if first_state_sram_input_id = 4177 then
	sram_write <= x"CC9C0010";
end if;
if first_state_sram_input_id = 4178 then
	sram_write <= x"CC7C0018";
end if;
if first_state_sram_input_id = 4179 then
	sram_write <= x"CCDC0020";
end if;
if first_state_sram_input_id = 4180 then
	sram_write <= x"C43C0028";
end if;
if first_state_sram_input_id = 4181 then
	sram_write <= x"CC5C0030";
end if;
if first_state_sram_input_id = 4182 then
	sram_write <= x"CCBC0038";
end if;
if first_state_sram_input_id = 4183 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 4184 then
	sram_write <= x"4020C000";
end if;
if first_state_sram_input_id = 4185 then
	sram_write <= x"03DC0048";
end if;
if first_state_sram_input_id = 4186 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 4187 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 4188 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 4189 then
	sram_write <= x"07DC0048";
end if;
if first_state_sram_input_id = 4190 then
	sram_write <= x"C85C0038";
end if;
if first_state_sram_input_id = 4191 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 4192 then
	sram_write <= x"C85C0030";
end if;
if first_state_sram_input_id = 4193 then
	sram_write <= x"44242000";
end if;
if first_state_sram_input_id = 4194 then
	sram_write <= x"C03C0028";
end if;
if first_state_sram_input_id = 4195 then
	sram_write <= x"CC220004";
end if;
if first_state_sram_input_id = 4196 then
	sram_write <= x"C05C0004";
end if;
if first_state_sram_input_id = 4197 then
	sram_write <= x"C8240008";
end if;
if first_state_sram_input_id = 4198 then
	sram_write <= x"C07C0000";
end if;
if first_state_sram_input_id = 4199 then
	sram_write <= x"C0860024";
end if;
if first_state_sram_input_id = 4200 then
	sram_write <= x"C8480000";
end if;
if first_state_sram_input_id = 4201 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 4202 then
	sram_write <= x"C8440000";
end if;
if first_state_sram_input_id = 4203 then
	sram_write <= x"C0860024";
end if;
if first_state_sram_input_id = 4204 then
	sram_write <= x"C8680008";
end if;
if first_state_sram_input_id = 4205 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 4206 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 4207 then
	sram_write <= x"C85C0020";
end if;
if first_state_sram_input_id = 4208 then
	sram_write <= x"CC3C0040";
end if;
if first_state_sram_input_id = 4209 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 4210 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 4211 then
	sram_write <= x"03DC0050";
end if;
if first_state_sram_input_id = 4212 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 4213 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 4214 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 4215 then
	sram_write <= x"07DC0050";
end if;
if first_state_sram_input_id = 4216 then
	sram_write <= x"C85C0040";
end if;
if first_state_sram_input_id = 4217 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 4218 then
	sram_write <= x"C85C0018";
end if;
if first_state_sram_input_id = 4219 then
	sram_write <= x"44242000";
end if;
if first_state_sram_input_id = 4220 then
	sram_write <= x"C03C0028";
end if;
if first_state_sram_input_id = 4221 then
	sram_write <= x"CC220008";
end if;
if first_state_sram_input_id = 4222 then
	sram_write <= x"C05C0004";
end if;
if first_state_sram_input_id = 4223 then
	sram_write <= x"C8240004";
end if;
if first_state_sram_input_id = 4224 then
	sram_write <= x"C07C0000";
end if;
if first_state_sram_input_id = 4225 then
	sram_write <= x"C0860024";
end if;
if first_state_sram_input_id = 4226 then
	sram_write <= x"C8480000";
end if;
if first_state_sram_input_id = 4227 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 4228 then
	sram_write <= x"C8440000";
end if;
if first_state_sram_input_id = 4229 then
	sram_write <= x"C0460024";
end if;
if first_state_sram_input_id = 4230 then
	sram_write <= x"C8640004";
end if;
if first_state_sram_input_id = 4231 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 4232 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 4233 then
	sram_write <= x"C85C0020";
end if;
if first_state_sram_input_id = 4234 then
	sram_write <= x"CC3C0048";
end if;
if first_state_sram_input_id = 4235 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 4236 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 4237 then
	sram_write <= x"03DC0058";
end if;
if first_state_sram_input_id = 4238 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 4239 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 4240 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 4241 then
	sram_write <= x"07DC0058";
end if;
if first_state_sram_input_id = 4242 then
	sram_write <= x"C85C0048";
end if;
if first_state_sram_input_id = 4243 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 4244 then
	sram_write <= x"C85C0010";
end if;
if first_state_sram_input_id = 4245 then
	sram_write <= x"44242000";
end if;
if first_state_sram_input_id = 4246 then
	sram_write <= x"C03C0028";
end if;
if first_state_sram_input_id = 4247 then
	sram_write <= x"CC22000C";
end if;
if first_state_sram_input_id = 4248 then
	sram_write <= x"82004270";
end if;
if first_state_sram_input_id = 4249 then
	sram_write <= x"CC420004";
end if;
if first_state_sram_input_id = 4250 then
	sram_write <= x"CC620008";
end if;
if first_state_sram_input_id = 4251 then
	sram_write <= x"CC82000C";
end if;
if first_state_sram_input_id = 4252 then
	sram_write <= x"C83C0008";
end if;
if first_state_sram_input_id = 4253 then
	sram_write <= x"8A2042A0";
end if;
if first_state_sram_input_id = 4254 then
	sram_write <= x"C43C0028";
end if;
if first_state_sram_input_id = 4255 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 4256 then
	sram_write <= x"03DC0058";
end if;
if first_state_sram_input_id = 4257 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 4258 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 4259 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 4260 then
	sram_write <= x"07DC0058";
end if;
if first_state_sram_input_id = 4261 then
	sram_write <= x"C03C0028";
end if;
if first_state_sram_input_id = 4262 then
	sram_write <= x"CC220010";
end if;
if first_state_sram_input_id = 4263 then
	sram_write <= x"820042A0";
end if;
if first_state_sram_input_id = 4264 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 4265 then
	sram_write <= x"86404628";
end if;
if first_state_sram_input_id = 4266 then
	sram_write <= x"026000C8";
end if;
if first_state_sram_input_id = 4267 then
	sram_write <= x"22840220";
end if;
if first_state_sram_input_id = 4268 then
	sram_write <= x"D0868000";
end if;
if first_state_sram_input_id = 4269 then
	sram_write <= x"C0A20004";
end if;
if first_state_sram_input_id = 4270 then
	sram_write <= x"C0C20000";
end if;
if first_state_sram_input_id = 4271 then
	sram_write <= x"C0E80004";
end if;
if first_state_sram_input_id = 4272 then
	sram_write <= x"03000001";
end if;
if first_state_sram_input_id = 4273 then
	sram_write <= x"C43C0000";
end if;
if first_state_sram_input_id = 4274 then
	sram_write <= x"C47C0004";
end if;
if first_state_sram_input_id = 4275 then
	sram_write <= x"82F04350";
end if;
if first_state_sram_input_id = 4276 then
	sram_write <= x"03000002";
end if;
if first_state_sram_input_id = 4277 then
	sram_write <= x"82F04314";
end if;
if first_state_sram_input_id = 4278 then
	sram_write <= x"C4BC0008";
end if;
if first_state_sram_input_id = 4279 then
	sram_write <= x"C45C000C";
end if;
if first_state_sram_input_id = 4280 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 4281 then
	sram_write <= x"00480000";
end if;
if first_state_sram_input_id = 4282 then
	sram_write <= x"002C0000";
end if;
if first_state_sram_input_id = 4283 then
	sram_write <= x"03DC0018";
end if;
if first_state_sram_input_id = 4284 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 4285 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 4286 then
	sram_write <= x"8200400C";
end if;
if first_state_sram_input_id = 4287 then
	sram_write <= x"07DC0018";
end if;
if first_state_sram_input_id = 4288 then
	sram_write <= x"C05C000C";
end if;
if first_state_sram_input_id = 4289 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 4290 then
	sram_write <= x"C09C0008";
end if;
if first_state_sram_input_id = 4291 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 4292 then
	sram_write <= x"8200434C";
end if;
if first_state_sram_input_id = 4293 then
	sram_write <= x"C4BC0008";
end if;
if first_state_sram_input_id = 4294 then
	sram_write <= x"C45C000C";
end if;
if first_state_sram_input_id = 4295 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 4296 then
	sram_write <= x"00480000";
end if;
if first_state_sram_input_id = 4297 then
	sram_write <= x"002C0000";
end if;
if first_state_sram_input_id = 4298 then
	sram_write <= x"03DC0018";
end if;
if first_state_sram_input_id = 4299 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 4300 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 4301 then
	sram_write <= x"82003E98";
end if;
if first_state_sram_input_id = 4302 then
	sram_write <= x"07DC0018";
end if;
if first_state_sram_input_id = 4303 then
	sram_write <= x"C05C000C";
end if;
if first_state_sram_input_id = 4304 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 4305 then
	sram_write <= x"C09C0008";
end if;
if first_state_sram_input_id = 4306 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 4307 then
	sram_write <= x"82004388";
end if;
if first_state_sram_input_id = 4308 then
	sram_write <= x"C4BC0008";
end if;
if first_state_sram_input_id = 4309 then
	sram_write <= x"C45C000C";
end if;
if first_state_sram_input_id = 4310 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 4311 then
	sram_write <= x"00480000";
end if;
if first_state_sram_input_id = 4312 then
	sram_write <= x"002C0000";
end if;
if first_state_sram_input_id = 4313 then
	sram_write <= x"03DC0018";
end if;
if first_state_sram_input_id = 4314 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 4315 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 4316 then
	sram_write <= x"82003CC4";
end if;
if first_state_sram_input_id = 4317 then
	sram_write <= x"07DC0018";
end if;
if first_state_sram_input_id = 4318 then
	sram_write <= x"C05C000C";
end if;
if first_state_sram_input_id = 4319 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 4320 then
	sram_write <= x"C09C0008";
end if;
if first_state_sram_input_id = 4321 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 4322 then
	sram_write <= x"06240001";
end if;
if first_state_sram_input_id = 4323 then
	sram_write <= x"86204624";
end if;
if first_state_sram_input_id = 4324 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 4325 then
	sram_write <= x"C07C0004";
end if;
if first_state_sram_input_id = 4326 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 4327 then
	sram_write <= x"C09C0000";
end if;
if first_state_sram_input_id = 4328 then
	sram_write <= x"C0A80004";
end if;
if first_state_sram_input_id = 4329 then
	sram_write <= x"C0C80000";
end if;
if first_state_sram_input_id = 4330 then
	sram_write <= x"C0E40004";
end if;
if first_state_sram_input_id = 4331 then
	sram_write <= x"03000001";
end if;
if first_state_sram_input_id = 4332 then
	sram_write <= x"82F0442C";
end if;
if first_state_sram_input_id = 4333 then
	sram_write <= x"03000002";
end if;
if first_state_sram_input_id = 4334 then
	sram_write <= x"82F043F4";
end if;
if first_state_sram_input_id = 4335 then
	sram_write <= x"C4BC0010";
end if;
if first_state_sram_input_id = 4336 then
	sram_write <= x"C43C0014";
end if;
if first_state_sram_input_id = 4337 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 4338 then
	sram_write <= x"002C0000";
end if;
if first_state_sram_input_id = 4339 then
	sram_write <= x"03DC0020";
end if;
if first_state_sram_input_id = 4340 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 4341 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 4342 then
	sram_write <= x"8200400C";
end if;
if first_state_sram_input_id = 4343 then
	sram_write <= x"07DC0020";
end if;
if first_state_sram_input_id = 4344 then
	sram_write <= x"C05C0014";
end if;
if first_state_sram_input_id = 4345 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 4346 then
	sram_write <= x"C09C0010";
end if;
if first_state_sram_input_id = 4347 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 4348 then
	sram_write <= x"82004428";
end if;
if first_state_sram_input_id = 4349 then
	sram_write <= x"C4BC0010";
end if;
if first_state_sram_input_id = 4350 then
	sram_write <= x"C43C0014";
end if;
if first_state_sram_input_id = 4351 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 4352 then
	sram_write <= x"002C0000";
end if;
if first_state_sram_input_id = 4353 then
	sram_write <= x"03DC0020";
end if;
if first_state_sram_input_id = 4354 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 4355 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 4356 then
	sram_write <= x"82003E98";
end if;
if first_state_sram_input_id = 4357 then
	sram_write <= x"07DC0020";
end if;
if first_state_sram_input_id = 4358 then
	sram_write <= x"C05C0014";
end if;
if first_state_sram_input_id = 4359 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 4360 then
	sram_write <= x"C09C0010";
end if;
if first_state_sram_input_id = 4361 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 4362 then
	sram_write <= x"82004460";
end if;
if first_state_sram_input_id = 4363 then
	sram_write <= x"C4BC0010";
end if;
if first_state_sram_input_id = 4364 then
	sram_write <= x"C43C0014";
end if;
if first_state_sram_input_id = 4365 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 4366 then
	sram_write <= x"002C0000";
end if;
if first_state_sram_input_id = 4367 then
	sram_write <= x"03DC0020";
end if;
if first_state_sram_input_id = 4368 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 4369 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 4370 then
	sram_write <= x"82003CC4";
end if;
if first_state_sram_input_id = 4371 then
	sram_write <= x"07DC0020";
end if;
if first_state_sram_input_id = 4372 then
	sram_write <= x"C05C0014";
end if;
if first_state_sram_input_id = 4373 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 4374 then
	sram_write <= x"C09C0010";
end if;
if first_state_sram_input_id = 4375 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 4376 then
	sram_write <= x"06240001";
end if;
if first_state_sram_input_id = 4377 then
	sram_write <= x"86204620";
end if;
if first_state_sram_input_id = 4378 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 4379 then
	sram_write <= x"C07C0004";
end if;
if first_state_sram_input_id = 4380 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 4381 then
	sram_write <= x"C09C0000";
end if;
if first_state_sram_input_id = 4382 then
	sram_write <= x"C0A80004";
end if;
if first_state_sram_input_id = 4383 then
	sram_write <= x"C0C80000";
end if;
if first_state_sram_input_id = 4384 then
	sram_write <= x"C0E40004";
end if;
if first_state_sram_input_id = 4385 then
	sram_write <= x"03000001";
end if;
if first_state_sram_input_id = 4386 then
	sram_write <= x"82F04504";
end if;
if first_state_sram_input_id = 4387 then
	sram_write <= x"03000002";
end if;
if first_state_sram_input_id = 4388 then
	sram_write <= x"82F044CC";
end if;
if first_state_sram_input_id = 4389 then
	sram_write <= x"C4BC0018";
end if;
if first_state_sram_input_id = 4390 then
	sram_write <= x"C43C001C";
end if;
if first_state_sram_input_id = 4391 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 4392 then
	sram_write <= x"002C0000";
end if;
if first_state_sram_input_id = 4393 then
	sram_write <= x"03DC0028";
end if;
if first_state_sram_input_id = 4394 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 4395 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 4396 then
	sram_write <= x"8200400C";
end if;
if first_state_sram_input_id = 4397 then
	sram_write <= x"07DC0028";
end if;
if first_state_sram_input_id = 4398 then
	sram_write <= x"C05C001C";
end if;
if first_state_sram_input_id = 4399 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 4400 then
	sram_write <= x"C09C0018";
end if;
if first_state_sram_input_id = 4401 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 4402 then
	sram_write <= x"82004500";
end if;
if first_state_sram_input_id = 4403 then
	sram_write <= x"C4BC0018";
end if;
if first_state_sram_input_id = 4404 then
	sram_write <= x"C43C001C";
end if;
if first_state_sram_input_id = 4405 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 4406 then
	sram_write <= x"002C0000";
end if;
if first_state_sram_input_id = 4407 then
	sram_write <= x"03DC0028";
end if;
if first_state_sram_input_id = 4408 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 4409 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 4410 then
	sram_write <= x"82003E98";
end if;
if first_state_sram_input_id = 4411 then
	sram_write <= x"07DC0028";
end if;
if first_state_sram_input_id = 4412 then
	sram_write <= x"C05C001C";
end if;
if first_state_sram_input_id = 4413 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 4414 then
	sram_write <= x"C09C0018";
end if;
if first_state_sram_input_id = 4415 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 4416 then
	sram_write <= x"82004538";
end if;
if first_state_sram_input_id = 4417 then
	sram_write <= x"C4BC0018";
end if;
if first_state_sram_input_id = 4418 then
	sram_write <= x"C43C001C";
end if;
if first_state_sram_input_id = 4419 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 4420 then
	sram_write <= x"002C0000";
end if;
if first_state_sram_input_id = 4421 then
	sram_write <= x"03DC0028";
end if;
if first_state_sram_input_id = 4422 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 4423 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 4424 then
	sram_write <= x"82003CC4";
end if;
if first_state_sram_input_id = 4425 then
	sram_write <= x"07DC0028";
end if;
if first_state_sram_input_id = 4426 then
	sram_write <= x"C05C001C";
end if;
if first_state_sram_input_id = 4427 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 4428 then
	sram_write <= x"C09C0018";
end if;
if first_state_sram_input_id = 4429 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 4430 then
	sram_write <= x"06240001";
end if;
if first_state_sram_input_id = 4431 then
	sram_write <= x"8620461C";
end if;
if first_state_sram_input_id = 4432 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 4433 then
	sram_write <= x"C07C0004";
end if;
if first_state_sram_input_id = 4434 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 4435 then
	sram_write <= x"C07C0000";
end if;
if first_state_sram_input_id = 4436 then
	sram_write <= x"C0860004";
end if;
if first_state_sram_input_id = 4437 then
	sram_write <= x"C0A60000";
end if;
if first_state_sram_input_id = 4438 then
	sram_write <= x"C0C40004";
end if;
if first_state_sram_input_id = 4439 then
	sram_write <= x"02E00001";
end if;
if first_state_sram_input_id = 4440 then
	sram_write <= x"82CE45DC";
end if;
if first_state_sram_input_id = 4441 then
	sram_write <= x"02E00002";
end if;
if first_state_sram_input_id = 4442 then
	sram_write <= x"82CE45A4";
end if;
if first_state_sram_input_id = 4443 then
	sram_write <= x"C49C0020";
end if;
if first_state_sram_input_id = 4444 then
	sram_write <= x"C43C0024";
end if;
if first_state_sram_input_id = 4445 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 4446 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 4447 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 4448 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 4449 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 4450 then
	sram_write <= x"8200400C";
end if;
if first_state_sram_input_id = 4451 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 4452 then
	sram_write <= x"C05C0024";
end if;
if first_state_sram_input_id = 4453 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 4454 then
	sram_write <= x"C09C0020";
end if;
if first_state_sram_input_id = 4455 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 4456 then
	sram_write <= x"820045D8";
end if;
if first_state_sram_input_id = 4457 then
	sram_write <= x"C49C0020";
end if;
if first_state_sram_input_id = 4458 then
	sram_write <= x"C43C0024";
end if;
if first_state_sram_input_id = 4459 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 4460 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 4461 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 4462 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 4463 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 4464 then
	sram_write <= x"82003E98";
end if;
if first_state_sram_input_id = 4465 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 4466 then
	sram_write <= x"C05C0024";
end if;
if first_state_sram_input_id = 4467 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 4468 then
	sram_write <= x"C09C0020";
end if;
if first_state_sram_input_id = 4469 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 4470 then
	sram_write <= x"82004610";
end if;
if first_state_sram_input_id = 4471 then
	sram_write <= x"C49C0020";
end if;
if first_state_sram_input_id = 4472 then
	sram_write <= x"C43C0024";
end if;
if first_state_sram_input_id = 4473 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 4474 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 4475 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 4476 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 4477 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 4478 then
	sram_write <= x"82003CC4";
end if;
if first_state_sram_input_id = 4479 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 4480 then
	sram_write <= x"C05C0024";
end if;
if first_state_sram_input_id = 4481 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 4482 then
	sram_write <= x"C09C0020";
end if;
if first_state_sram_input_id = 4483 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 4484 then
	sram_write <= x"06440001";
end if;
if first_state_sram_input_id = 4485 then
	sram_write <= x"C03C0000";
end if;
if first_state_sram_input_id = 4486 then
	sram_write <= x"820042A4";
end if;
if first_state_sram_input_id = 4487 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 4488 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 4489 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 4490 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 4491 then
	sram_write <= x"8640477C";
end if;
if first_state_sram_input_id = 4492 then
	sram_write <= x"026000C8";
end if;
if first_state_sram_input_id = 4493 then
	sram_write <= x"22840220";
end if;
if first_state_sram_input_id = 4494 then
	sram_write <= x"D0668000";
end if;
if first_state_sram_input_id = 4495 then
	sram_write <= x"C0860028";
end if;
if first_state_sram_input_id = 4496 then
	sram_write <= x"C0A60004";
end if;
if first_state_sram_input_id = 4497 then
	sram_write <= x"C8220000";
end if;
if first_state_sram_input_id = 4498 then
	sram_write <= x"C0C60014";
end if;
if first_state_sram_input_id = 4499 then
	sram_write <= x"C84C0000";
end if;
if first_state_sram_input_id = 4500 then
	sram_write <= x"44224000";
end if;
if first_state_sram_input_id = 4501 then
	sram_write <= x"CC280000";
end if;
if first_state_sram_input_id = 4502 then
	sram_write <= x"C8220004";
end if;
if first_state_sram_input_id = 4503 then
	sram_write <= x"C0C60014";
end if;
if first_state_sram_input_id = 4504 then
	sram_write <= x"C84C0004";
end if;
if first_state_sram_input_id = 4505 then
	sram_write <= x"44224000";
end if;
if first_state_sram_input_id = 4506 then
	sram_write <= x"CC280004";
end if;
if first_state_sram_input_id = 4507 then
	sram_write <= x"C8220008";
end if;
if first_state_sram_input_id = 4508 then
	sram_write <= x"C0C60014";
end if;
if first_state_sram_input_id = 4509 then
	sram_write <= x"C84C0008";
end if;
if first_state_sram_input_id = 4510 then
	sram_write <= x"44224000";
end if;
if first_state_sram_input_id = 4511 then
	sram_write <= x"CC280008";
end if;
if first_state_sram_input_id = 4512 then
	sram_write <= x"02C00002";
end if;
if first_state_sram_input_id = 4513 then
	sram_write <= x"82AC4740";
end if;
if first_state_sram_input_id = 4514 then
	sram_write <= x"02C00002";
end if;
if first_state_sram_input_id = 4515 then
	sram_write <= x"86CA4694";
end if;
if first_state_sram_input_id = 4516 then
	sram_write <= x"8200473C";
end if;
if first_state_sram_input_id = 4517 then
	sram_write <= x"C8280000";
end if;
if first_state_sram_input_id = 4518 then
	sram_write <= x"C8480004";
end if;
if first_state_sram_input_id = 4519 then
	sram_write <= x"C8680008";
end if;
if first_state_sram_input_id = 4520 then
	sram_write <= x"48822000";
end if;
if first_state_sram_input_id = 4521 then
	sram_write <= x"C0C60010";
end if;
if first_state_sram_input_id = 4522 then
	sram_write <= x"C8AC0000";
end if;
if first_state_sram_input_id = 4523 then
	sram_write <= x"4888A000";
end if;
if first_state_sram_input_id = 4524 then
	sram_write <= x"48A44000";
end if;
if first_state_sram_input_id = 4525 then
	sram_write <= x"C0C60010";
end if;
if first_state_sram_input_id = 4526 then
	sram_write <= x"C8CC0004";
end if;
if first_state_sram_input_id = 4527 then
	sram_write <= x"48AAC000";
end if;
if first_state_sram_input_id = 4528 then
	sram_write <= x"4088A000";
end if;
if first_state_sram_input_id = 4529 then
	sram_write <= x"48A66000";
end if;
if first_state_sram_input_id = 4530 then
	sram_write <= x"C0C60010";
end if;
if first_state_sram_input_id = 4531 then
	sram_write <= x"C8CC0008";
end if;
if first_state_sram_input_id = 4532 then
	sram_write <= x"48AAC000";
end if;
if first_state_sram_input_id = 4533 then
	sram_write <= x"4088A000";
end if;
if first_state_sram_input_id = 4534 then
	sram_write <= x"C0C6000C";
end if;
if first_state_sram_input_id = 4535 then
	sram_write <= x"82C04720";
end if;
if first_state_sram_input_id = 4536 then
	sram_write <= x"48A46000";
end if;
if first_state_sram_input_id = 4537 then
	sram_write <= x"C0C60024";
end if;
if first_state_sram_input_id = 4538 then
	sram_write <= x"C8CC0000";
end if;
if first_state_sram_input_id = 4539 then
	sram_write <= x"48AAC000";
end if;
if first_state_sram_input_id = 4540 then
	sram_write <= x"4088A000";
end if;
if first_state_sram_input_id = 4541 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 4542 then
	sram_write <= x"C0C60024";
end if;
if first_state_sram_input_id = 4543 then
	sram_write <= x"C8AC0004";
end if;
if first_state_sram_input_id = 4544 then
	sram_write <= x"4866A000";
end if;
if first_state_sram_input_id = 4545 then
	sram_write <= x"40686000";
end if;
if first_state_sram_input_id = 4546 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 4547 then
	sram_write <= x"C0660024";
end if;
if first_state_sram_input_id = 4548 then
	sram_write <= x"C8460008";
end if;
if first_state_sram_input_id = 4549 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 4550 then
	sram_write <= x"40262000";
end if;
if first_state_sram_input_id = 4551 then
	sram_write <= x"82004724";
end if;
if first_state_sram_input_id = 4552 then
	sram_write <= x"40208000";
end if;
if first_state_sram_input_id = 4553 then
	sram_write <= x"02600003";
end if;
if first_state_sram_input_id = 4554 then
	sram_write <= x"82A64730";
end if;
if first_state_sram_input_id = 4555 then
	sram_write <= x"82004738";
end if;
if first_state_sram_input_id = 4556 then
	sram_write <= x"C84000A8";
end if;
if first_state_sram_input_id = 4557 then
	sram_write <= x"44224000";
end if;
if first_state_sram_input_id = 4558 then
	sram_write <= x"CC28000C";
end if;
if first_state_sram_input_id = 4559 then
	sram_write <= x"82004774";
end if;
if first_state_sram_input_id = 4560 then
	sram_write <= x"C0660010";
end if;
if first_state_sram_input_id = 4561 then
	sram_write <= x"C8280000";
end if;
if first_state_sram_input_id = 4562 then
	sram_write <= x"C8480004";
end if;
if first_state_sram_input_id = 4563 then
	sram_write <= x"C8680008";
end if;
if first_state_sram_input_id = 4564 then
	sram_write <= x"C8860000";
end if;
if first_state_sram_input_id = 4565 then
	sram_write <= x"48282000";
end if;
if first_state_sram_input_id = 4566 then
	sram_write <= x"C8860004";
end if;
if first_state_sram_input_id = 4567 then
	sram_write <= x"48484000";
end if;
if first_state_sram_input_id = 4568 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 4569 then
	sram_write <= x"C8460008";
end if;
if first_state_sram_input_id = 4570 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 4571 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 4572 then
	sram_write <= x"CC28000C";
end if;
if first_state_sram_input_id = 4573 then
	sram_write <= x"06440001";
end if;
if first_state_sram_input_id = 4574 then
	sram_write <= x"8200462C";
end if;
if first_state_sram_input_id = 4575 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 4576 then
	sram_write <= x"48822000";
end if;
if first_state_sram_input_id = 4577 then
	sram_write <= x"C0420010";
end if;
if first_state_sram_input_id = 4578 then
	sram_write <= x"C8A40000";
end if;
if first_state_sram_input_id = 4579 then
	sram_write <= x"4888A000";
end if;
if first_state_sram_input_id = 4580 then
	sram_write <= x"48A44000";
end if;
if first_state_sram_input_id = 4581 then
	sram_write <= x"C0420010";
end if;
if first_state_sram_input_id = 4582 then
	sram_write <= x"C8C40004";
end if;
if first_state_sram_input_id = 4583 then
	sram_write <= x"48AAC000";
end if;
if first_state_sram_input_id = 4584 then
	sram_write <= x"4088A000";
end if;
if first_state_sram_input_id = 4585 then
	sram_write <= x"48A66000";
end if;
if first_state_sram_input_id = 4586 then
	sram_write <= x"C0420010";
end if;
if first_state_sram_input_id = 4587 then
	sram_write <= x"C8C40008";
end if;
if first_state_sram_input_id = 4588 then
	sram_write <= x"48AAC000";
end if;
if first_state_sram_input_id = 4589 then
	sram_write <= x"4088A000";
end if;
if first_state_sram_input_id = 4590 then
	sram_write <= x"C042000C";
end if;
if first_state_sram_input_id = 4591 then
	sram_write <= x"82404800";
end if;
if first_state_sram_input_id = 4592 then
	sram_write <= x"48A46000";
end if;
if first_state_sram_input_id = 4593 then
	sram_write <= x"C0420024";
end if;
if first_state_sram_input_id = 4594 then
	sram_write <= x"C8C40000";
end if;
if first_state_sram_input_id = 4595 then
	sram_write <= x"48AAC000";
end if;
if first_state_sram_input_id = 4596 then
	sram_write <= x"4088A000";
end if;
if first_state_sram_input_id = 4597 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 4598 then
	sram_write <= x"C0420024";
end if;
if first_state_sram_input_id = 4599 then
	sram_write <= x"C8A40004";
end if;
if first_state_sram_input_id = 4600 then
	sram_write <= x"4866A000";
end if;
if first_state_sram_input_id = 4601 then
	sram_write <= x"40686000";
end if;
if first_state_sram_input_id = 4602 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 4603 then
	sram_write <= x"C0420024";
end if;
if first_state_sram_input_id = 4604 then
	sram_write <= x"C8440008";
end if;
if first_state_sram_input_id = 4605 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 4606 then
	sram_write <= x"40262000";
end if;
if first_state_sram_input_id = 4607 then
	sram_write <= x"82004804";
end if;
if first_state_sram_input_id = 4608 then
	sram_write <= x"40208000";
end if;
if first_state_sram_input_id = 4609 then
	sram_write <= x"C0420004";
end if;
if first_state_sram_input_id = 4610 then
	sram_write <= x"02600003";
end if;
if first_state_sram_input_id = 4611 then
	sram_write <= x"82464814";
end if;
if first_state_sram_input_id = 4612 then
	sram_write <= x"8200481C";
end if;
if first_state_sram_input_id = 4613 then
	sram_write <= x"C84000A8";
end if;
if first_state_sram_input_id = 4614 then
	sram_write <= x"44224000";
end if;
if first_state_sram_input_id = 4615 then
	sram_write <= x"C0220018";
end if;
if first_state_sram_input_id = 4616 then
	sram_write <= x"8E20482C";
end if;
if first_state_sram_input_id = 4617 then
	sram_write <= x"02400000";
end if;
if first_state_sram_input_id = 4618 then
	sram_write <= x"82004830";
end if;
if first_state_sram_input_id = 4619 then
	sram_write <= x"02400001";
end if;
if first_state_sram_input_id = 4620 then
	sram_write <= x"82204848";
end if;
if first_state_sram_input_id = 4621 then
	sram_write <= x"8E204840";
end if;
if first_state_sram_input_id = 4622 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 4623 then
	sram_write <= x"82004844";
end if;
if first_state_sram_input_id = 4624 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 4625 then
	sram_write <= x"8200484C";
end if;
if first_state_sram_input_id = 4626 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 4627 then
	sram_write <= x"82204858";
end if;
if first_state_sram_input_id = 4628 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 4629 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 4630 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 4631 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 4632 then
	sram_write <= x"C0420014";
end if;
if first_state_sram_input_id = 4633 then
	sram_write <= x"C8840000";
end if;
if first_state_sram_input_id = 4634 then
	sram_write <= x"44228000";
end if;
if first_state_sram_input_id = 4635 then
	sram_write <= x"C0420014";
end if;
if first_state_sram_input_id = 4636 then
	sram_write <= x"C8840004";
end if;
if first_state_sram_input_id = 4637 then
	sram_write <= x"44448000";
end if;
if first_state_sram_input_id = 4638 then
	sram_write <= x"C0420014";
end if;
if first_state_sram_input_id = 4639 then
	sram_write <= x"C8840008";
end if;
if first_state_sram_input_id = 4640 then
	sram_write <= x"44668000";
end if;
if first_state_sram_input_id = 4641 then
	sram_write <= x"C0420004";
end if;
if first_state_sram_input_id = 4642 then
	sram_write <= x"02600001";
end if;
if first_state_sram_input_id = 4643 then
	sram_write <= x"8246497C";
end if;
if first_state_sram_input_id = 4644 then
	sram_write <= x"02600002";
end if;
if first_state_sram_input_id = 4645 then
	sram_write <= x"82464914";
end if;
if first_state_sram_input_id = 4646 then
	sram_write <= x"C43C0000";
end if;
if first_state_sram_input_id = 4647 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 4648 then
	sram_write <= x"03DC000C";
end if;
if first_state_sram_input_id = 4649 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 4650 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 4651 then
	sram_write <= x"82003344";
end if;
if first_state_sram_input_id = 4652 then
	sram_write <= x"07DC000C";
end if;
if first_state_sram_input_id = 4653 then
	sram_write <= x"C03C0000";
end if;
if first_state_sram_input_id = 4654 then
	sram_write <= x"C0420004";
end if;
if first_state_sram_input_id = 4655 then
	sram_write <= x"02600003";
end if;
if first_state_sram_input_id = 4656 then
	sram_write <= x"824648C8";
end if;
if first_state_sram_input_id = 4657 then
	sram_write <= x"820048D0";
end if;
if first_state_sram_input_id = 4658 then
	sram_write <= x"C84000A8";
end if;
if first_state_sram_input_id = 4659 then
	sram_write <= x"44224000";
end if;
if first_state_sram_input_id = 4660 then
	sram_write <= x"C0220018";
end if;
if first_state_sram_input_id = 4661 then
	sram_write <= x"8E2048E0";
end if;
if first_state_sram_input_id = 4662 then
	sram_write <= x"02400000";
end if;
if first_state_sram_input_id = 4663 then
	sram_write <= x"820048E4";
end if;
if first_state_sram_input_id = 4664 then
	sram_write <= x"02400001";
end if;
if first_state_sram_input_id = 4665 then
	sram_write <= x"822048FC";
end if;
if first_state_sram_input_id = 4666 then
	sram_write <= x"8E2048F4";
end if;
if first_state_sram_input_id = 4667 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 4668 then
	sram_write <= x"820048F8";
end if;
if first_state_sram_input_id = 4669 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 4670 then
	sram_write <= x"82004900";
end if;
if first_state_sram_input_id = 4671 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 4672 then
	sram_write <= x"8220490C";
end if;
if first_state_sram_input_id = 4673 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 4674 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 4675 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 4676 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 4677 then
	sram_write <= x"C0420010";
end if;
if first_state_sram_input_id = 4678 then
	sram_write <= x"C8840000";
end if;
if first_state_sram_input_id = 4679 then
	sram_write <= x"48282000";
end if;
if first_state_sram_input_id = 4680 then
	sram_write <= x"C8840004";
end if;
if first_state_sram_input_id = 4681 then
	sram_write <= x"48484000";
end if;
if first_state_sram_input_id = 4682 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 4683 then
	sram_write <= x"C8440008";
end if;
if first_state_sram_input_id = 4684 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 4685 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 4686 then
	sram_write <= x"C0220018";
end if;
if first_state_sram_input_id = 4687 then
	sram_write <= x"8E204948";
end if;
if first_state_sram_input_id = 4688 then
	sram_write <= x"02400000";
end if;
if first_state_sram_input_id = 4689 then
	sram_write <= x"8200494C";
end if;
if first_state_sram_input_id = 4690 then
	sram_write <= x"02400001";
end if;
if first_state_sram_input_id = 4691 then
	sram_write <= x"82204964";
end if;
if first_state_sram_input_id = 4692 then
	sram_write <= x"8E20495C";
end if;
if first_state_sram_input_id = 4693 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 4694 then
	sram_write <= x"82004960";
end if;
if first_state_sram_input_id = 4695 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 4696 then
	sram_write <= x"82004968";
end if;
if first_state_sram_input_id = 4697 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 4698 then
	sram_write <= x"82204974";
end if;
if first_state_sram_input_id = 4699 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 4700 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 4701 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 4702 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 4703 then
	sram_write <= x"8E204984";
end if;
if first_state_sram_input_id = 4704 then
	sram_write <= x"82004988";
end if;
if first_state_sram_input_id = 4705 then
	sram_write <= x"44202000";
end if;
if first_state_sram_input_id = 4706 then
	sram_write <= x"C0420010";
end if;
if first_state_sram_input_id = 4707 then
	sram_write <= x"C8840000";
end if;
if first_state_sram_input_id = 4708 then
	sram_write <= x"8E28499C";
end if;
if first_state_sram_input_id = 4709 then
	sram_write <= x"02400000";
end if;
if first_state_sram_input_id = 4710 then
	sram_write <= x"820049E8";
end if;
if first_state_sram_input_id = 4711 then
	sram_write <= x"8E4049A8";
end if;
if first_state_sram_input_id = 4712 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 4713 then
	sram_write <= x"820049AC";
end if;
if first_state_sram_input_id = 4714 then
	sram_write <= x"44204000";
end if;
if first_state_sram_input_id = 4715 then
	sram_write <= x"C0420010";
end if;
if first_state_sram_input_id = 4716 then
	sram_write <= x"C8440004";
end if;
if first_state_sram_input_id = 4717 then
	sram_write <= x"8E2449C0";
end if;
if first_state_sram_input_id = 4718 then
	sram_write <= x"02400000";
end if;
if first_state_sram_input_id = 4719 then
	sram_write <= x"820049E8";
end if;
if first_state_sram_input_id = 4720 then
	sram_write <= x"8E6049CC";
end if;
if first_state_sram_input_id = 4721 then
	sram_write <= x"40206000";
end if;
if first_state_sram_input_id = 4722 then
	sram_write <= x"820049D0";
end if;
if first_state_sram_input_id = 4723 then
	sram_write <= x"44206000";
end if;
if first_state_sram_input_id = 4724 then
	sram_write <= x"C0420010";
end if;
if first_state_sram_input_id = 4725 then
	sram_write <= x"C8440008";
end if;
if first_state_sram_input_id = 4726 then
	sram_write <= x"8E2449E4";
end if;
if first_state_sram_input_id = 4727 then
	sram_write <= x"02400000";
end if;
if first_state_sram_input_id = 4728 then
	sram_write <= x"820049E8";
end if;
if first_state_sram_input_id = 4729 then
	sram_write <= x"02400001";
end if;
if first_state_sram_input_id = 4730 then
	sram_write <= x"824049F4";
end if;
if first_state_sram_input_id = 4731 then
	sram_write <= x"C0220018";
end if;
if first_state_sram_input_id = 4732 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 4733 then
	sram_write <= x"C0220018";
end if;
if first_state_sram_input_id = 4734 then
	sram_write <= x"82204A04";
end if;
if first_state_sram_input_id = 4735 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 4736 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 4737 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 4738 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 4739 then
	sram_write <= x"22620220";
end if;
if first_state_sram_input_id = 4740 then
	sram_write <= x"D0646000";
end if;
if first_state_sram_input_id = 4741 then
	sram_write <= x"0280FFFF";
end if;
if first_state_sram_input_id = 4742 then
	sram_write <= x"82684E38";
end if;
if first_state_sram_input_id = 4743 then
	sram_write <= x"028000C8";
end if;
if first_state_sram_input_id = 4744 then
	sram_write <= x"22660220";
end if;
if first_state_sram_input_id = 4745 then
	sram_write <= x"D0686000";
end if;
if first_state_sram_input_id = 4746 then
	sram_write <= x"C0A60014";
end if;
if first_state_sram_input_id = 4747 then
	sram_write <= x"C88A0000";
end if;
if first_state_sram_input_id = 4748 then
	sram_write <= x"44828000";
end if;
if first_state_sram_input_id = 4749 then
	sram_write <= x"C0A60014";
end if;
if first_state_sram_input_id = 4750 then
	sram_write <= x"C8AA0004";
end if;
if first_state_sram_input_id = 4751 then
	sram_write <= x"44A4A000";
end if;
if first_state_sram_input_id = 4752 then
	sram_write <= x"C0A60014";
end if;
if first_state_sram_input_id = 4753 then
	sram_write <= x"C8CA0008";
end if;
if first_state_sram_input_id = 4754 then
	sram_write <= x"44C6C000";
end if;
if first_state_sram_input_id = 4755 then
	sram_write <= x"C0A60004";
end if;
if first_state_sram_input_id = 4756 then
	sram_write <= x"02C00001";
end if;
if first_state_sram_input_id = 4757 then
	sram_write <= x"CC7C0000";
end if;
if first_state_sram_input_id = 4758 then
	sram_write <= x"CC5C0008";
end if;
if first_state_sram_input_id = 4759 then
	sram_write <= x"CC3C0010";
end if;
if first_state_sram_input_id = 4760 then
	sram_write <= x"C49C0018";
end if;
if first_state_sram_input_id = 4761 then
	sram_write <= x"C45C001C";
end if;
if first_state_sram_input_id = 4762 then
	sram_write <= x"C43C0020";
end if;
if first_state_sram_input_id = 4763 then
	sram_write <= x"82AC4B0C";
end if;
if first_state_sram_input_id = 4764 then
	sram_write <= x"02C00002";
end if;
if first_state_sram_input_id = 4765 then
	sram_write <= x"82AC4AA4";
end if;
if first_state_sram_input_id = 4766 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 4767 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 4768 then
	sram_write <= x"4060C000";
end if;
if first_state_sram_input_id = 4769 then
	sram_write <= x"4040A000";
end if;
if first_state_sram_input_id = 4770 then
	sram_write <= x"40208000";
end if;
if first_state_sram_input_id = 4771 then
	sram_write <= x"03DC002C";
end if;
if first_state_sram_input_id = 4772 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 4773 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 4774 then
	sram_write <= x"82004780";
end if;
if first_state_sram_input_id = 4775 then
	sram_write <= x"07DC002C";
end if;
if first_state_sram_input_id = 4776 then
	sram_write <= x"82004B08";
end if;
if first_state_sram_input_id = 4777 then
	sram_write <= x"C0A60010";
end if;
if first_state_sram_input_id = 4778 then
	sram_write <= x"C8EA0000";
end if;
if first_state_sram_input_id = 4779 then
	sram_write <= x"488E8000";
end if;
if first_state_sram_input_id = 4780 then
	sram_write <= x"C8EA0004";
end if;
if first_state_sram_input_id = 4781 then
	sram_write <= x"48AEA000";
end if;
if first_state_sram_input_id = 4782 then
	sram_write <= x"4088A000";
end if;
if first_state_sram_input_id = 4783 then
	sram_write <= x"C8AA0008";
end if;
if first_state_sram_input_id = 4784 then
	sram_write <= x"48AAC000";
end if;
if first_state_sram_input_id = 4785 then
	sram_write <= x"4088A000";
end if;
if first_state_sram_input_id = 4786 then
	sram_write <= x"C0660018";
end if;
if first_state_sram_input_id = 4787 then
	sram_write <= x"8E804AD8";
end if;
if first_state_sram_input_id = 4788 then
	sram_write <= x"02A00000";
end if;
if first_state_sram_input_id = 4789 then
	sram_write <= x"82004ADC";
end if;
if first_state_sram_input_id = 4790 then
	sram_write <= x"02A00001";
end if;
if first_state_sram_input_id = 4791 then
	sram_write <= x"82604AF4";
end if;
if first_state_sram_input_id = 4792 then
	sram_write <= x"8E804AEC";
end if;
if first_state_sram_input_id = 4793 then
	sram_write <= x"02600001";
end if;
if first_state_sram_input_id = 4794 then
	sram_write <= x"82004AF0";
end if;
if first_state_sram_input_id = 4795 then
	sram_write <= x"02600000";
end if;
if first_state_sram_input_id = 4796 then
	sram_write <= x"82004AF8";
end if;
if first_state_sram_input_id = 4797 then
	sram_write <= x"006A0000";
end if;
if first_state_sram_input_id = 4798 then
	sram_write <= x"82604B04";
end if;
if first_state_sram_input_id = 4799 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 4800 then
	sram_write <= x"82004B08";
end if;
if first_state_sram_input_id = 4801 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 4802 then
	sram_write <= x"82004B9C";
end if;
if first_state_sram_input_id = 4803 then
	sram_write <= x"8E804B14";
end if;
if first_state_sram_input_id = 4804 then
	sram_write <= x"82004B18";
end if;
if first_state_sram_input_id = 4805 then
	sram_write <= x"44808000";
end if;
if first_state_sram_input_id = 4806 then
	sram_write <= x"C0A60010";
end if;
if first_state_sram_input_id = 4807 then
	sram_write <= x"C8EA0000";
end if;
if first_state_sram_input_id = 4808 then
	sram_write <= x"8E8E4B2C";
end if;
if first_state_sram_input_id = 4809 then
	sram_write <= x"02A00000";
end if;
if first_state_sram_input_id = 4810 then
	sram_write <= x"82004B78";
end if;
if first_state_sram_input_id = 4811 then
	sram_write <= x"8EA04B38";
end if;
if first_state_sram_input_id = 4812 then
	sram_write <= x"4080A000";
end if;
if first_state_sram_input_id = 4813 then
	sram_write <= x"82004B3C";
end if;
if first_state_sram_input_id = 4814 then
	sram_write <= x"4480A000";
end if;
if first_state_sram_input_id = 4815 then
	sram_write <= x"C0A60010";
end if;
if first_state_sram_input_id = 4816 then
	sram_write <= x"C8AA0004";
end if;
if first_state_sram_input_id = 4817 then
	sram_write <= x"8E8A4B50";
end if;
if first_state_sram_input_id = 4818 then
	sram_write <= x"02A00000";
end if;
if first_state_sram_input_id = 4819 then
	sram_write <= x"82004B78";
end if;
if first_state_sram_input_id = 4820 then
	sram_write <= x"8EC04B5C";
end if;
if first_state_sram_input_id = 4821 then
	sram_write <= x"4080C000";
end if;
if first_state_sram_input_id = 4822 then
	sram_write <= x"82004B60";
end if;
if first_state_sram_input_id = 4823 then
	sram_write <= x"4480C000";
end if;
if first_state_sram_input_id = 4824 then
	sram_write <= x"C0A60010";
end if;
if first_state_sram_input_id = 4825 then
	sram_write <= x"C8AA0008";
end if;
if first_state_sram_input_id = 4826 then
	sram_write <= x"8E8A4B74";
end if;
if first_state_sram_input_id = 4827 then
	sram_write <= x"02A00000";
end if;
if first_state_sram_input_id = 4828 then
	sram_write <= x"82004B78";
end if;
if first_state_sram_input_id = 4829 then
	sram_write <= x"02A00001";
end if;
if first_state_sram_input_id = 4830 then
	sram_write <= x"82A04B88";
end if;
if first_state_sram_input_id = 4831 then
	sram_write <= x"C0660018";
end if;
if first_state_sram_input_id = 4832 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 4833 then
	sram_write <= x"82004B9C";
end if;
if first_state_sram_input_id = 4834 then
	sram_write <= x"C0660018";
end if;
if first_state_sram_input_id = 4835 then
	sram_write <= x"82604B98";
end if;
if first_state_sram_input_id = 4836 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 4837 then
	sram_write <= x"82004B9C";
end if;
if first_state_sram_input_id = 4838 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 4839 then
	sram_write <= x"82204BA8";
end if;
if first_state_sram_input_id = 4840 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 4841 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 4842 then
	sram_write <= x"C03C0020";
end if;
if first_state_sram_input_id = 4843 then
	sram_write <= x"02220001";
end if;
if first_state_sram_input_id = 4844 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 4845 then
	sram_write <= x"C07C001C";
end if;
if first_state_sram_input_id = 4846 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 4847 then
	sram_write <= x"0280FFFF";
end if;
if first_state_sram_input_id = 4848 then
	sram_write <= x"82484E30";
end if;
if first_state_sram_input_id = 4849 then
	sram_write <= x"22440220";
end if;
if first_state_sram_input_id = 4850 then
	sram_write <= x"C09C0018";
end if;
if first_state_sram_input_id = 4851 then
	sram_write <= x"D0484000";
end if;
if first_state_sram_input_id = 4852 then
	sram_write <= x"C83C0010";
end if;
if first_state_sram_input_id = 4853 then
	sram_write <= x"C85C0008";
end if;
if first_state_sram_input_id = 4854 then
	sram_write <= x"C87C0000";
end if;
if first_state_sram_input_id = 4855 then
	sram_write <= x"C43C0024";
end if;
if first_state_sram_input_id = 4856 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 4857 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 4858 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 4859 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 4860 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 4861 then
	sram_write <= x"82004860";
end if;
if first_state_sram_input_id = 4862 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 4863 then
	sram_write <= x"82204C08";
end if;
if first_state_sram_input_id = 4864 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 4865 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 4866 then
	sram_write <= x"C03C0024";
end if;
if first_state_sram_input_id = 4867 then
	sram_write <= x"02220001";
end if;
if first_state_sram_input_id = 4868 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 4869 then
	sram_write <= x"C07C001C";
end if;
if first_state_sram_input_id = 4870 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 4871 then
	sram_write <= x"0280FFFF";
end if;
if first_state_sram_input_id = 4872 then
	sram_write <= x"82484E28";
end if;
if first_state_sram_input_id = 4873 then
	sram_write <= x"22440220";
end if;
if first_state_sram_input_id = 4874 then
	sram_write <= x"C09C0018";
end if;
if first_state_sram_input_id = 4875 then
	sram_write <= x"D0484000";
end if;
if first_state_sram_input_id = 4876 then
	sram_write <= x"C0A40014";
end if;
if first_state_sram_input_id = 4877 then
	sram_write <= x"C82A0000";
end if;
if first_state_sram_input_id = 4878 then
	sram_write <= x"C85C0010";
end if;
if first_state_sram_input_id = 4879 then
	sram_write <= x"44242000";
end if;
if first_state_sram_input_id = 4880 then
	sram_write <= x"C0A40014";
end if;
if first_state_sram_input_id = 4881 then
	sram_write <= x"C86A0004";
end if;
if first_state_sram_input_id = 4882 then
	sram_write <= x"C89C0008";
end if;
if first_state_sram_input_id = 4883 then
	sram_write <= x"44686000";
end if;
if first_state_sram_input_id = 4884 then
	sram_write <= x"C0A40014";
end if;
if first_state_sram_input_id = 4885 then
	sram_write <= x"C8AA0008";
end if;
if first_state_sram_input_id = 4886 then
	sram_write <= x"C8DC0000";
end if;
if first_state_sram_input_id = 4887 then
	sram_write <= x"44ACA000";
end if;
if first_state_sram_input_id = 4888 then
	sram_write <= x"C0A40004";
end if;
if first_state_sram_input_id = 4889 then
	sram_write <= x"02C00001";
end if;
if first_state_sram_input_id = 4890 then
	sram_write <= x"C43C0028";
end if;
if first_state_sram_input_id = 4891 then
	sram_write <= x"82AC4D08";
end if;
if first_state_sram_input_id = 4892 then
	sram_write <= x"02C00002";
end if;
if first_state_sram_input_id = 4893 then
	sram_write <= x"82AC4CA0";
end if;
if first_state_sram_input_id = 4894 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 4895 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 4896 then
	sram_write <= x"40406000";
end if;
if first_state_sram_input_id = 4897 then
	sram_write <= x"4060A000";
end if;
if first_state_sram_input_id = 4898 then
	sram_write <= x"03DC0034";
end if;
if first_state_sram_input_id = 4899 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 4900 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 4901 then
	sram_write <= x"82004780";
end if;
if first_state_sram_input_id = 4902 then
	sram_write <= x"07DC0034";
end if;
if first_state_sram_input_id = 4903 then
	sram_write <= x"82004D04";
end if;
if first_state_sram_input_id = 4904 then
	sram_write <= x"C0A40010";
end if;
if first_state_sram_input_id = 4905 then
	sram_write <= x"C8EA0000";
end if;
if first_state_sram_input_id = 4906 then
	sram_write <= x"482E2000";
end if;
if first_state_sram_input_id = 4907 then
	sram_write <= x"C8EA0004";
end if;
if first_state_sram_input_id = 4908 then
	sram_write <= x"486E6000";
end if;
if first_state_sram_input_id = 4909 then
	sram_write <= x"40226000";
end if;
if first_state_sram_input_id = 4910 then
	sram_write <= x"C86A0008";
end if;
if first_state_sram_input_id = 4911 then
	sram_write <= x"4866A000";
end if;
if first_state_sram_input_id = 4912 then
	sram_write <= x"40226000";
end if;
if first_state_sram_input_id = 4913 then
	sram_write <= x"C0440018";
end if;
if first_state_sram_input_id = 4914 then
	sram_write <= x"8E204CD4";
end if;
if first_state_sram_input_id = 4915 then
	sram_write <= x"02A00000";
end if;
if first_state_sram_input_id = 4916 then
	sram_write <= x"82004CD8";
end if;
if first_state_sram_input_id = 4917 then
	sram_write <= x"02A00001";
end if;
if first_state_sram_input_id = 4918 then
	sram_write <= x"82404CF0";
end if;
if first_state_sram_input_id = 4919 then
	sram_write <= x"8E204CE8";
end if;
if first_state_sram_input_id = 4920 then
	sram_write <= x"02400001";
end if;
if first_state_sram_input_id = 4921 then
	sram_write <= x"82004CEC";
end if;
if first_state_sram_input_id = 4922 then
	sram_write <= x"02400000";
end if;
if first_state_sram_input_id = 4923 then
	sram_write <= x"82004CF4";
end if;
if first_state_sram_input_id = 4924 then
	sram_write <= x"004A0000";
end if;
if first_state_sram_input_id = 4925 then
	sram_write <= x"82404D00";
end if;
if first_state_sram_input_id = 4926 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 4927 then
	sram_write <= x"82004D04";
end if;
if first_state_sram_input_id = 4928 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 4929 then
	sram_write <= x"82004D98";
end if;
if first_state_sram_input_id = 4930 then
	sram_write <= x"8E204D10";
end if;
if first_state_sram_input_id = 4931 then
	sram_write <= x"82004D14";
end if;
if first_state_sram_input_id = 4932 then
	sram_write <= x"44202000";
end if;
if first_state_sram_input_id = 4933 then
	sram_write <= x"C0A40010";
end if;
if first_state_sram_input_id = 4934 then
	sram_write <= x"C8EA0000";
end if;
if first_state_sram_input_id = 4935 then
	sram_write <= x"8E2E4D28";
end if;
if first_state_sram_input_id = 4936 then
	sram_write <= x"02A00000";
end if;
if first_state_sram_input_id = 4937 then
	sram_write <= x"82004D74";
end if;
if first_state_sram_input_id = 4938 then
	sram_write <= x"8E604D34";
end if;
if first_state_sram_input_id = 4939 then
	sram_write <= x"40206000";
end if;
if first_state_sram_input_id = 4940 then
	sram_write <= x"82004D38";
end if;
if first_state_sram_input_id = 4941 then
	sram_write <= x"44206000";
end if;
if first_state_sram_input_id = 4942 then
	sram_write <= x"C0A40010";
end if;
if first_state_sram_input_id = 4943 then
	sram_write <= x"C86A0004";
end if;
if first_state_sram_input_id = 4944 then
	sram_write <= x"8E264D4C";
end if;
if first_state_sram_input_id = 4945 then
	sram_write <= x"02A00000";
end if;
if first_state_sram_input_id = 4946 then
	sram_write <= x"82004D74";
end if;
if first_state_sram_input_id = 4947 then
	sram_write <= x"8EA04D58";
end if;
if first_state_sram_input_id = 4948 then
	sram_write <= x"4020A000";
end if;
if first_state_sram_input_id = 4949 then
	sram_write <= x"82004D5C";
end if;
if first_state_sram_input_id = 4950 then
	sram_write <= x"4420A000";
end if;
if first_state_sram_input_id = 4951 then
	sram_write <= x"C0A40010";
end if;
if first_state_sram_input_id = 4952 then
	sram_write <= x"C86A0008";
end if;
if first_state_sram_input_id = 4953 then
	sram_write <= x"8E264D70";
end if;
if first_state_sram_input_id = 4954 then
	sram_write <= x"02A00000";
end if;
if first_state_sram_input_id = 4955 then
	sram_write <= x"82004D74";
end if;
if first_state_sram_input_id = 4956 then
	sram_write <= x"02A00001";
end if;
if first_state_sram_input_id = 4957 then
	sram_write <= x"82A04D84";
end if;
if first_state_sram_input_id = 4958 then
	sram_write <= x"C0440018";
end if;
if first_state_sram_input_id = 4959 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 4960 then
	sram_write <= x"82004D98";
end if;
if first_state_sram_input_id = 4961 then
	sram_write <= x"C0440018";
end if;
if first_state_sram_input_id = 4962 then
	sram_write <= x"82404D94";
end if;
if first_state_sram_input_id = 4963 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 4964 then
	sram_write <= x"82004D98";
end if;
if first_state_sram_input_id = 4965 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 4966 then
	sram_write <= x"82204DA4";
end if;
if first_state_sram_input_id = 4967 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 4968 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 4969 then
	sram_write <= x"C03C0028";
end if;
if first_state_sram_input_id = 4970 then
	sram_write <= x"02220001";
end if;
if first_state_sram_input_id = 4971 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 4972 then
	sram_write <= x"C07C001C";
end if;
if first_state_sram_input_id = 4973 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 4974 then
	sram_write <= x"0280FFFF";
end if;
if first_state_sram_input_id = 4975 then
	sram_write <= x"82484E20";
end if;
if first_state_sram_input_id = 4976 then
	sram_write <= x"22440220";
end if;
if first_state_sram_input_id = 4977 then
	sram_write <= x"C09C0018";
end if;
if first_state_sram_input_id = 4978 then
	sram_write <= x"D0484000";
end if;
if first_state_sram_input_id = 4979 then
	sram_write <= x"C83C0010";
end if;
if first_state_sram_input_id = 4980 then
	sram_write <= x"C85C0008";
end if;
if first_state_sram_input_id = 4981 then
	sram_write <= x"C87C0000";
end if;
if first_state_sram_input_id = 4982 then
	sram_write <= x"C43C002C";
end if;
if first_state_sram_input_id = 4983 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 4984 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 4985 then
	sram_write <= x"03DC0038";
end if;
if first_state_sram_input_id = 4986 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 4987 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 4988 then
	sram_write <= x"82004860";
end if;
if first_state_sram_input_id = 4989 then
	sram_write <= x"07DC0038";
end if;
if first_state_sram_input_id = 4990 then
	sram_write <= x"82204E04";
end if;
if first_state_sram_input_id = 4991 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 4992 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 4993 then
	sram_write <= x"C03C002C";
end if;
if first_state_sram_input_id = 4994 then
	sram_write <= x"02220001";
end if;
if first_state_sram_input_id = 4995 then
	sram_write <= x"C83C0010";
end if;
if first_state_sram_input_id = 4996 then
	sram_write <= x"C85C0008";
end if;
if first_state_sram_input_id = 4997 then
	sram_write <= x"C87C0000";
end if;
if first_state_sram_input_id = 4998 then
	sram_write <= x"C05C001C";
end if;
if first_state_sram_input_id = 4999 then
	sram_write <= x"82004A0C";
end if;
if first_state_sram_input_id = 5000 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 5001 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 5002 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 5003 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 5004 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 5005 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 5006 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 5007 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 5008 then
	sram_write <= x"22620220";
end if;
if first_state_sram_input_id = 5009 then
	sram_write <= x"D0646000";
end if;
if first_state_sram_input_id = 5010 then
	sram_write <= x"0280FFFF";
end if;
if first_state_sram_input_id = 5011 then
	sram_write <= x"8268527C";
end if;
if first_state_sram_input_id = 5012 then
	sram_write <= x"02800368";
end if;
if first_state_sram_input_id = 5013 then
	sram_write <= x"02A002B8";
end if;
if first_state_sram_input_id = 5014 then
	sram_write <= x"02C000C8";
end if;
if first_state_sram_input_id = 5015 then
	sram_write <= x"22E60220";
end if;
if first_state_sram_input_id = 5016 then
	sram_write <= x"D0ECE000";
end if;
if first_state_sram_input_id = 5017 then
	sram_write <= x"C82A0000";
end if;
if first_state_sram_input_id = 5018 then
	sram_write <= x"C10E0014";
end if;
if first_state_sram_input_id = 5019 then
	sram_write <= x"C8500000";
end if;
if first_state_sram_input_id = 5020 then
	sram_write <= x"44224000";
end if;
if first_state_sram_input_id = 5021 then
	sram_write <= x"C84A0004";
end if;
if first_state_sram_input_id = 5022 then
	sram_write <= x"C10E0014";
end if;
if first_state_sram_input_id = 5023 then
	sram_write <= x"C8700004";
end if;
if first_state_sram_input_id = 5024 then
	sram_write <= x"44446000";
end if;
if first_state_sram_input_id = 5025 then
	sram_write <= x"C86A0008";
end if;
if first_state_sram_input_id = 5026 then
	sram_write <= x"C10E0014";
end if;
if first_state_sram_input_id = 5027 then
	sram_write <= x"C8900008";
end if;
if first_state_sram_input_id = 5028 then
	sram_write <= x"44668000";
end if;
if first_state_sram_input_id = 5029 then
	sram_write <= x"C1080004";
end if;
if first_state_sram_input_id = 5030 then
	sram_write <= x"23260220";
end if;
if first_state_sram_input_id = 5031 then
	sram_write <= x"D1112000";
end if;
if first_state_sram_input_id = 5032 then
	sram_write <= x"C12E0004";
end if;
if first_state_sram_input_id = 5033 then
	sram_write <= x"03400001";
end if;
if first_state_sram_input_id = 5034 then
	sram_write <= x"C4BC0000";
end if;
if first_state_sram_input_id = 5035 then
	sram_write <= x"C45C0004";
end if;
if first_state_sram_input_id = 5036 then
	sram_write <= x"C43C0008";
end if;
if first_state_sram_input_id = 5037 then
	sram_write <= x"C4DC000C";
end if;
if first_state_sram_input_id = 5038 then
	sram_write <= x"C47C0010";
end if;
if first_state_sram_input_id = 5039 then
	sram_write <= x"83344F2C";
end if;
if first_state_sram_input_id = 5040 then
	sram_write <= x"02800002";
end if;
if first_state_sram_input_id = 5041 then
	sram_write <= x"83284EEC";
end if;
if first_state_sram_input_id = 5042 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 5043 then
	sram_write <= x"00500000";
end if;
if first_state_sram_input_id = 5044 then
	sram_write <= x"002E0000";
end if;
if first_state_sram_input_id = 5045 then
	sram_write <= x"03DC001C";
end if;
if first_state_sram_input_id = 5046 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 5047 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 5048 then
	sram_write <= x"82003A54";
end if;
if first_state_sram_input_id = 5049 then
	sram_write <= x"07DC001C";
end if;
if first_state_sram_input_id = 5050 then
	sram_write <= x"82004F28";
end if;
if first_state_sram_input_id = 5051 then
	sram_write <= x"C8900000";
end if;
if first_state_sram_input_id = 5052 then
	sram_write <= x"8E804EFC";
end if;
if first_state_sram_input_id = 5053 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 5054 then
	sram_write <= x"82004F28";
end if;
if first_state_sram_input_id = 5055 then
	sram_write <= x"028002AC";
end if;
if first_state_sram_input_id = 5056 then
	sram_write <= x"C8900004";
end if;
if first_state_sram_input_id = 5057 then
	sram_write <= x"48282000";
end if;
if first_state_sram_input_id = 5058 then
	sram_write <= x"C8900008";
end if;
if first_state_sram_input_id = 5059 then
	sram_write <= x"48484000";
end if;
if first_state_sram_input_id = 5060 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 5061 then
	sram_write <= x"C850000C";
end if;
if first_state_sram_input_id = 5062 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 5063 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 5064 then
	sram_write <= x"CC280000";
end if;
if first_state_sram_input_id = 5065 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 5066 then
	sram_write <= x"82004F54";
end if;
if first_state_sram_input_id = 5067 then
	sram_write <= x"C0880000";
end if;
if first_state_sram_input_id = 5068 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 5069 then
	sram_write <= x"00700000";
end if;
if first_state_sram_input_id = 5070 then
	sram_write <= x"00480000";
end if;
if first_state_sram_input_id = 5071 then
	sram_write <= x"002E0000";
end if;
if first_state_sram_input_id = 5072 then
	sram_write <= x"03DC001C";
end if;
if first_state_sram_input_id = 5073 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 5074 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 5075 then
	sram_write <= x"8200389C";
end if;
if first_state_sram_input_id = 5076 then
	sram_write <= x"07DC001C";
end if;
if first_state_sram_input_id = 5077 then
	sram_write <= x"024002AC";
end if;
if first_state_sram_input_id = 5078 then
	sram_write <= x"C8240000";
end if;
if first_state_sram_input_id = 5079 then
	sram_write <= x"82204F78";
end if;
if first_state_sram_input_id = 5080 then
	sram_write <= x"C8400078";
end if;
if first_state_sram_input_id = 5081 then
	sram_write <= x"8E244F70";
end if;
if first_state_sram_input_id = 5082 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 5083 then
	sram_write <= x"82004F74";
end if;
if first_state_sram_input_id = 5084 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 5085 then
	sram_write <= x"82004F7C";
end if;
if first_state_sram_input_id = 5086 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 5087 then
	sram_write <= x"8220524C";
end if;
if first_state_sram_input_id = 5088 then
	sram_write <= x"C8400074";
end if;
if first_state_sram_input_id = 5089 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 5090 then
	sram_write <= x"022001D0";
end if;
if first_state_sram_input_id = 5091 then
	sram_write <= x"C8420000";
end if;
if first_state_sram_input_id = 5092 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 5093 then
	sram_write <= x"C05C0000";
end if;
if first_state_sram_input_id = 5094 then
	sram_write <= x"C8640000";
end if;
if first_state_sram_input_id = 5095 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 5096 then
	sram_write <= x"C8620004";
end if;
if first_state_sram_input_id = 5097 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 5098 then
	sram_write <= x"C8840004";
end if;
if first_state_sram_input_id = 5099 then
	sram_write <= x"40668000";
end if;
if first_state_sram_input_id = 5100 then
	sram_write <= x"C8820008";
end if;
if first_state_sram_input_id = 5101 then
	sram_write <= x"48282000";
end if;
if first_state_sram_input_id = 5102 then
	sram_write <= x"C8840008";
end if;
if first_state_sram_input_id = 5103 then
	sram_write <= x"40228000";
end if;
if first_state_sram_input_id = 5104 then
	sram_write <= x"C05C0004";
end if;
if first_state_sram_input_id = 5105 then
	sram_write <= x"C0240000";
end if;
if first_state_sram_input_id = 5106 then
	sram_write <= x"0260FFFF";
end if;
if first_state_sram_input_id = 5107 then
	sram_write <= x"8226522C";
end if;
if first_state_sram_input_id = 5108 then
	sram_write <= x"22220220";
end if;
if first_state_sram_input_id = 5109 then
	sram_write <= x"C07C000C";
end if;
if first_state_sram_input_id = 5110 then
	sram_write <= x"D0262000";
end if;
if first_state_sram_input_id = 5111 then
	sram_write <= x"CC3C0018";
end if;
if first_state_sram_input_id = 5112 then
	sram_write <= x"CC7C0020";
end if;
if first_state_sram_input_id = 5113 then
	sram_write <= x"CC5C0028";
end if;
if first_state_sram_input_id = 5114 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 5115 then
	sram_write <= x"41E06000";
end if;
if first_state_sram_input_id = 5116 then
	sram_write <= x"40602000";
end if;
if first_state_sram_input_id = 5117 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 5118 then
	sram_write <= x"4041E000";
end if;
if first_state_sram_input_id = 5119 then
	sram_write <= x"03DC0038";
end if;
if first_state_sram_input_id = 5120 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 5121 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 5122 then
	sram_write <= x"82004860";
end if;
if first_state_sram_input_id = 5123 then
	sram_write <= x"07DC0038";
end if;
if first_state_sram_input_id = 5124 then
	sram_write <= x"8220501C";
end if;
if first_state_sram_input_id = 5125 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 5126 then
	sram_write <= x"82005228";
end if;
if first_state_sram_input_id = 5127 then
	sram_write <= x"C05C0004";
end if;
if first_state_sram_input_id = 5128 then
	sram_write <= x"C0240004";
end if;
if first_state_sram_input_id = 5129 then
	sram_write <= x"0260FFFF";
end if;
if first_state_sram_input_id = 5130 then
	sram_write <= x"82265224";
end if;
if first_state_sram_input_id = 5131 then
	sram_write <= x"22220220";
end if;
if first_state_sram_input_id = 5132 then
	sram_write <= x"C07C000C";
end if;
if first_state_sram_input_id = 5133 then
	sram_write <= x"D0262000";
end if;
if first_state_sram_input_id = 5134 then
	sram_write <= x"C0820014";
end if;
if first_state_sram_input_id = 5135 then
	sram_write <= x"C8280000";
end if;
if first_state_sram_input_id = 5136 then
	sram_write <= x"C85C0028";
end if;
if first_state_sram_input_id = 5137 then
	sram_write <= x"44242000";
end if;
if first_state_sram_input_id = 5138 then
	sram_write <= x"C0820014";
end if;
if first_state_sram_input_id = 5139 then
	sram_write <= x"C8680004";
end if;
if first_state_sram_input_id = 5140 then
	sram_write <= x"C89C0020";
end if;
if first_state_sram_input_id = 5141 then
	sram_write <= x"44686000";
end if;
if first_state_sram_input_id = 5142 then
	sram_write <= x"C0820014";
end if;
if first_state_sram_input_id = 5143 then
	sram_write <= x"C8A80008";
end if;
if first_state_sram_input_id = 5144 then
	sram_write <= x"C8DC0018";
end if;
if first_state_sram_input_id = 5145 then
	sram_write <= x"44ACA000";
end if;
if first_state_sram_input_id = 5146 then
	sram_write <= x"C0820004";
end if;
if first_state_sram_input_id = 5147 then
	sram_write <= x"02A00001";
end if;
if first_state_sram_input_id = 5148 then
	sram_write <= x"828A5108";
end if;
if first_state_sram_input_id = 5149 then
	sram_write <= x"02A00002";
end if;
if first_state_sram_input_id = 5150 then
	sram_write <= x"828A50A0";
end if;
if first_state_sram_input_id = 5151 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 5152 then
	sram_write <= x"40406000";
end if;
if first_state_sram_input_id = 5153 then
	sram_write <= x"4060A000";
end if;
if first_state_sram_input_id = 5154 then
	sram_write <= x"03DC0038";
end if;
if first_state_sram_input_id = 5155 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 5156 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 5157 then
	sram_write <= x"82004780";
end if;
if first_state_sram_input_id = 5158 then
	sram_write <= x"07DC0038";
end if;
if first_state_sram_input_id = 5159 then
	sram_write <= x"82005104";
end if;
if first_state_sram_input_id = 5160 then
	sram_write <= x"C0820010";
end if;
if first_state_sram_input_id = 5161 then
	sram_write <= x"C8E80000";
end if;
if first_state_sram_input_id = 5162 then
	sram_write <= x"482E2000";
end if;
if first_state_sram_input_id = 5163 then
	sram_write <= x"C8E80004";
end if;
if first_state_sram_input_id = 5164 then
	sram_write <= x"486E6000";
end if;
if first_state_sram_input_id = 5165 then
	sram_write <= x"40226000";
end if;
if first_state_sram_input_id = 5166 then
	sram_write <= x"C8680008";
end if;
if first_state_sram_input_id = 5167 then
	sram_write <= x"4866A000";
end if;
if first_state_sram_input_id = 5168 then
	sram_write <= x"40226000";
end if;
if first_state_sram_input_id = 5169 then
	sram_write <= x"C0220018";
end if;
if first_state_sram_input_id = 5170 then
	sram_write <= x"8E2050D4";
end if;
if first_state_sram_input_id = 5171 then
	sram_write <= x"02800000";
end if;
if first_state_sram_input_id = 5172 then
	sram_write <= x"820050D8";
end if;
if first_state_sram_input_id = 5173 then
	sram_write <= x"02800001";
end if;
if first_state_sram_input_id = 5174 then
	sram_write <= x"822050F0";
end if;
if first_state_sram_input_id = 5175 then
	sram_write <= x"8E2050E8";
end if;
if first_state_sram_input_id = 5176 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 5177 then
	sram_write <= x"820050EC";
end if;
if first_state_sram_input_id = 5178 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 5179 then
	sram_write <= x"820050F4";
end if;
if first_state_sram_input_id = 5180 then
	sram_write <= x"00280000";
end if;
if first_state_sram_input_id = 5181 then
	sram_write <= x"82205100";
end if;
if first_state_sram_input_id = 5182 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 5183 then
	sram_write <= x"82005104";
end if;
if first_state_sram_input_id = 5184 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 5185 then
	sram_write <= x"82005194";
end if;
if first_state_sram_input_id = 5186 then
	sram_write <= x"8E205110";
end if;
if first_state_sram_input_id = 5187 then
	sram_write <= x"82005114";
end if;
if first_state_sram_input_id = 5188 then
	sram_write <= x"44202000";
end if;
if first_state_sram_input_id = 5189 then
	sram_write <= x"C0820010";
end if;
if first_state_sram_input_id = 5190 then
	sram_write <= x"C8E80000";
end if;
if first_state_sram_input_id = 5191 then
	sram_write <= x"8E2E5128";
end if;
if first_state_sram_input_id = 5192 then
	sram_write <= x"02800000";
end if;
if first_state_sram_input_id = 5193 then
	sram_write <= x"82005174";
end if;
if first_state_sram_input_id = 5194 then
	sram_write <= x"8E605134";
end if;
if first_state_sram_input_id = 5195 then
	sram_write <= x"40206000";
end if;
if first_state_sram_input_id = 5196 then
	sram_write <= x"82005138";
end if;
if first_state_sram_input_id = 5197 then
	sram_write <= x"44206000";
end if;
if first_state_sram_input_id = 5198 then
	sram_write <= x"C0820010";
end if;
if first_state_sram_input_id = 5199 then
	sram_write <= x"C8680004";
end if;
if first_state_sram_input_id = 5200 then
	sram_write <= x"8E26514C";
end if;
if first_state_sram_input_id = 5201 then
	sram_write <= x"02800000";
end if;
if first_state_sram_input_id = 5202 then
	sram_write <= x"82005174";
end if;
if first_state_sram_input_id = 5203 then
	sram_write <= x"8EA05158";
end if;
if first_state_sram_input_id = 5204 then
	sram_write <= x"4020A000";
end if;
if first_state_sram_input_id = 5205 then
	sram_write <= x"8200515C";
end if;
if first_state_sram_input_id = 5206 then
	sram_write <= x"4420A000";
end if;
if first_state_sram_input_id = 5207 then
	sram_write <= x"C0820010";
end if;
if first_state_sram_input_id = 5208 then
	sram_write <= x"C8680008";
end if;
if first_state_sram_input_id = 5209 then
	sram_write <= x"8E265170";
end if;
if first_state_sram_input_id = 5210 then
	sram_write <= x"02800000";
end if;
if first_state_sram_input_id = 5211 then
	sram_write <= x"82005174";
end if;
if first_state_sram_input_id = 5212 then
	sram_write <= x"02800001";
end if;
if first_state_sram_input_id = 5213 then
	sram_write <= x"82805180";
end if;
if first_state_sram_input_id = 5214 then
	sram_write <= x"C0220018";
end if;
if first_state_sram_input_id = 5215 then
	sram_write <= x"82005194";
end if;
if first_state_sram_input_id = 5216 then
	sram_write <= x"C0220018";
end if;
if first_state_sram_input_id = 5217 then
	sram_write <= x"82205190";
end if;
if first_state_sram_input_id = 5218 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 5219 then
	sram_write <= x"82005194";
end if;
if first_state_sram_input_id = 5220 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 5221 then
	sram_write <= x"822051A0";
end if;
if first_state_sram_input_id = 5222 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 5223 then
	sram_write <= x"82005220";
end if;
if first_state_sram_input_id = 5224 then
	sram_write <= x"C05C0004";
end if;
if first_state_sram_input_id = 5225 then
	sram_write <= x"C0240008";
end if;
if first_state_sram_input_id = 5226 then
	sram_write <= x"0260FFFF";
end if;
if first_state_sram_input_id = 5227 then
	sram_write <= x"8226521C";
end if;
if first_state_sram_input_id = 5228 then
	sram_write <= x"22220220";
end if;
if first_state_sram_input_id = 5229 then
	sram_write <= x"C07C000C";
end if;
if first_state_sram_input_id = 5230 then
	sram_write <= x"D0262000";
end if;
if first_state_sram_input_id = 5231 then
	sram_write <= x"C83C0028";
end if;
if first_state_sram_input_id = 5232 then
	sram_write <= x"C85C0020";
end if;
if first_state_sram_input_id = 5233 then
	sram_write <= x"C87C0018";
end if;
if first_state_sram_input_id = 5234 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 5235 then
	sram_write <= x"03DC0038";
end if;
if first_state_sram_input_id = 5236 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 5237 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 5238 then
	sram_write <= x"82004860";
end if;
if first_state_sram_input_id = 5239 then
	sram_write <= x"07DC0038";
end if;
if first_state_sram_input_id = 5240 then
	sram_write <= x"822051EC";
end if;
if first_state_sram_input_id = 5241 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 5242 then
	sram_write <= x"82005218";
end if;
if first_state_sram_input_id = 5243 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 5244 then
	sram_write <= x"C83C0028";
end if;
if first_state_sram_input_id = 5245 then
	sram_write <= x"C85C0020";
end if;
if first_state_sram_input_id = 5246 then
	sram_write <= x"C87C0018";
end if;
if first_state_sram_input_id = 5247 then
	sram_write <= x"C05C0004";
end if;
if first_state_sram_input_id = 5248 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 5249 then
	sram_write <= x"03DC0038";
end if;
if first_state_sram_input_id = 5250 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 5251 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 5252 then
	sram_write <= x"82004A0C";
end if;
if first_state_sram_input_id = 5253 then
	sram_write <= x"07DC0038";
end if;
if first_state_sram_input_id = 5254 then
	sram_write <= x"82005220";
end if;
if first_state_sram_input_id = 5255 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 5256 then
	sram_write <= x"82005228";
end if;
if first_state_sram_input_id = 5257 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 5258 then
	sram_write <= x"82005230";
end if;
if first_state_sram_input_id = 5259 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 5260 then
	sram_write <= x"8220523C";
end if;
if first_state_sram_input_id = 5261 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 5262 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 5263 then
	sram_write <= x"C03C0008";
end if;
if first_state_sram_input_id = 5264 then
	sram_write <= x"02220001";
end if;
if first_state_sram_input_id = 5265 then
	sram_write <= x"C05C0004";
end if;
if first_state_sram_input_id = 5266 then
	sram_write <= x"82004E40";
end if;
if first_state_sram_input_id = 5267 then
	sram_write <= x"C03C0010";
end if;
if first_state_sram_input_id = 5268 then
	sram_write <= x"22220220";
end if;
if first_state_sram_input_id = 5269 then
	sram_write <= x"C05C000C";
end if;
if first_state_sram_input_id = 5270 then
	sram_write <= x"D0242000";
end if;
if first_state_sram_input_id = 5271 then
	sram_write <= x"C0220018";
end if;
if first_state_sram_input_id = 5272 then
	sram_write <= x"82205274";
end if;
if first_state_sram_input_id = 5273 then
	sram_write <= x"C03C0008";
end if;
if first_state_sram_input_id = 5274 then
	sram_write <= x"02220001";
end if;
if first_state_sram_input_id = 5275 then
	sram_write <= x"C05C0004";
end if;
if first_state_sram_input_id = 5276 then
	sram_write <= x"82004E40";
end if;
if first_state_sram_input_id = 5277 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 5278 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 5279 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 5280 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 5281 then
	sram_write <= x"22620220";
end if;
if first_state_sram_input_id = 5282 then
	sram_write <= x"D0646000";
end if;
if first_state_sram_input_id = 5283 then
	sram_write <= x"0280FFFF";
end if;
if first_state_sram_input_id = 5284 then
	sram_write <= x"8268540C";
end if;
if first_state_sram_input_id = 5285 then
	sram_write <= x"028001E0";
end if;
if first_state_sram_input_id = 5286 then
	sram_write <= x"22660220";
end if;
if first_state_sram_input_id = 5287 then
	sram_write <= x"D0686000";
end if;
if first_state_sram_input_id = 5288 then
	sram_write <= x"02A00000";
end if;
if first_state_sram_input_id = 5289 then
	sram_write <= x"C49C0000";
end if;
if first_state_sram_input_id = 5290 then
	sram_write <= x"C45C0004";
end if;
if first_state_sram_input_id = 5291 then
	sram_write <= x"C43C0008";
end if;
if first_state_sram_input_id = 5292 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 5293 then
	sram_write <= x"00460000";
end if;
if first_state_sram_input_id = 5294 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 5295 then
	sram_write <= x"03DC0014";
end if;
if first_state_sram_input_id = 5296 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 5297 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 5298 then
	sram_write <= x"82004E40";
end if;
if first_state_sram_input_id = 5299 then
	sram_write <= x"07DC0014";
end if;
if first_state_sram_input_id = 5300 then
	sram_write <= x"822052DC";
end if;
if first_state_sram_input_id = 5301 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 5302 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 5303 then
	sram_write <= x"C03C0008";
end if;
if first_state_sram_input_id = 5304 then
	sram_write <= x"02220001";
end if;
if first_state_sram_input_id = 5305 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 5306 then
	sram_write <= x"C07C0004";
end if;
if first_state_sram_input_id = 5307 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 5308 then
	sram_write <= x"0280FFFF";
end if;
if first_state_sram_input_id = 5309 then
	sram_write <= x"82485404";
end if;
if first_state_sram_input_id = 5310 then
	sram_write <= x"22440220";
end if;
if first_state_sram_input_id = 5311 then
	sram_write <= x"C09C0000";
end if;
if first_state_sram_input_id = 5312 then
	sram_write <= x"D0484000";
end if;
if first_state_sram_input_id = 5313 then
	sram_write <= x"02A00000";
end if;
if first_state_sram_input_id = 5314 then
	sram_write <= x"C43C000C";
end if;
if first_state_sram_input_id = 5315 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 5316 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 5317 then
	sram_write <= x"03DC0018";
end if;
if first_state_sram_input_id = 5318 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 5319 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 5320 then
	sram_write <= x"82004E40";
end if;
if first_state_sram_input_id = 5321 then
	sram_write <= x"07DC0018";
end if;
if first_state_sram_input_id = 5322 then
	sram_write <= x"82205334";
end if;
if first_state_sram_input_id = 5323 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 5324 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 5325 then
	sram_write <= x"C03C000C";
end if;
if first_state_sram_input_id = 5326 then
	sram_write <= x"02220001";
end if;
if first_state_sram_input_id = 5327 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 5328 then
	sram_write <= x"C07C0004";
end if;
if first_state_sram_input_id = 5329 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 5330 then
	sram_write <= x"0280FFFF";
end if;
if first_state_sram_input_id = 5331 then
	sram_write <= x"824853FC";
end if;
if first_state_sram_input_id = 5332 then
	sram_write <= x"22440220";
end if;
if first_state_sram_input_id = 5333 then
	sram_write <= x"C09C0000";
end if;
if first_state_sram_input_id = 5334 then
	sram_write <= x"D0484000";
end if;
if first_state_sram_input_id = 5335 then
	sram_write <= x"02A00000";
end if;
if first_state_sram_input_id = 5336 then
	sram_write <= x"C43C0010";
end if;
if first_state_sram_input_id = 5337 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 5338 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 5339 then
	sram_write <= x"03DC001C";
end if;
if first_state_sram_input_id = 5340 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 5341 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 5342 then
	sram_write <= x"82004E40";
end if;
if first_state_sram_input_id = 5343 then
	sram_write <= x"07DC001C";
end if;
if first_state_sram_input_id = 5344 then
	sram_write <= x"8220538C";
end if;
if first_state_sram_input_id = 5345 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 5346 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 5347 then
	sram_write <= x"C03C0010";
end if;
if first_state_sram_input_id = 5348 then
	sram_write <= x"02220001";
end if;
if first_state_sram_input_id = 5349 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 5350 then
	sram_write <= x"C07C0004";
end if;
if first_state_sram_input_id = 5351 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 5352 then
	sram_write <= x"0280FFFF";
end if;
if first_state_sram_input_id = 5353 then
	sram_write <= x"824853F4";
end if;
if first_state_sram_input_id = 5354 then
	sram_write <= x"22440220";
end if;
if first_state_sram_input_id = 5355 then
	sram_write <= x"C09C0000";
end if;
if first_state_sram_input_id = 5356 then
	sram_write <= x"D0484000";
end if;
if first_state_sram_input_id = 5357 then
	sram_write <= x"02800000";
end if;
if first_state_sram_input_id = 5358 then
	sram_write <= x"C43C0014";
end if;
if first_state_sram_input_id = 5359 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 5360 then
	sram_write <= x"00280000";
end if;
if first_state_sram_input_id = 5361 then
	sram_write <= x"03DC0020";
end if;
if first_state_sram_input_id = 5362 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 5363 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 5364 then
	sram_write <= x"82004E40";
end if;
if first_state_sram_input_id = 5365 then
	sram_write <= x"07DC0020";
end if;
if first_state_sram_input_id = 5366 then
	sram_write <= x"822053E4";
end if;
if first_state_sram_input_id = 5367 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 5368 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 5369 then
	sram_write <= x"C03C0014";
end if;
if first_state_sram_input_id = 5370 then
	sram_write <= x"02220001";
end if;
if first_state_sram_input_id = 5371 then
	sram_write <= x"C05C0004";
end if;
if first_state_sram_input_id = 5372 then
	sram_write <= x"82005284";
end if;
if first_state_sram_input_id = 5373 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 5374 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 5375 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 5376 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 5377 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 5378 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 5379 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 5380 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 5381 then
	sram_write <= x"22620220";
end if;
if first_state_sram_input_id = 5382 then
	sram_write <= x"D0646000";
end if;
if first_state_sram_input_id = 5383 then
	sram_write <= x"C0860000";
end if;
if first_state_sram_input_id = 5384 then
	sram_write <= x"02A0FFFF";
end if;
if first_state_sram_input_id = 5385 then
	sram_write <= x"828A57C0";
end if;
if first_state_sram_input_id = 5386 then
	sram_write <= x"02A00063";
end if;
if first_state_sram_input_id = 5387 then
	sram_write <= x"C47C0000";
end if;
if first_state_sram_input_id = 5388 then
	sram_write <= x"C45C0004";
end if;
if first_state_sram_input_id = 5389 then
	sram_write <= x"C43C0008";
end if;
if first_state_sram_input_id = 5390 then
	sram_write <= x"828A5678";
end if;
if first_state_sram_input_id = 5391 then
	sram_write <= x"02A00368";
end if;
if first_state_sram_input_id = 5392 then
	sram_write <= x"02C002B8";
end if;
if first_state_sram_input_id = 5393 then
	sram_write <= x"02E000C8";
end if;
if first_state_sram_input_id = 5394 then
	sram_write <= x"23080220";
end if;
if first_state_sram_input_id = 5395 then
	sram_write <= x"D0EF0000";
end if;
if first_state_sram_input_id = 5396 then
	sram_write <= x"C82C0000";
end if;
if first_state_sram_input_id = 5397 then
	sram_write <= x"C10E0014";
end if;
if first_state_sram_input_id = 5398 then
	sram_write <= x"C8500000";
end if;
if first_state_sram_input_id = 5399 then
	sram_write <= x"44224000";
end if;
if first_state_sram_input_id = 5400 then
	sram_write <= x"C84C0004";
end if;
if first_state_sram_input_id = 5401 then
	sram_write <= x"C10E0014";
end if;
if first_state_sram_input_id = 5402 then
	sram_write <= x"C8700004";
end if;
if first_state_sram_input_id = 5403 then
	sram_write <= x"44446000";
end if;
if first_state_sram_input_id = 5404 then
	sram_write <= x"C86C0008";
end if;
if first_state_sram_input_id = 5405 then
	sram_write <= x"C0CE0014";
end if;
if first_state_sram_input_id = 5406 then
	sram_write <= x"C88C0008";
end if;
if first_state_sram_input_id = 5407 then
	sram_write <= x"44668000";
end if;
if first_state_sram_input_id = 5408 then
	sram_write <= x"C0CA0004";
end if;
if first_state_sram_input_id = 5409 then
	sram_write <= x"22880220";
end if;
if first_state_sram_input_id = 5410 then
	sram_write <= x"D08C8000";
end if;
if first_state_sram_input_id = 5411 then
	sram_write <= x"C0CE0004";
end if;
if first_state_sram_input_id = 5412 then
	sram_write <= x"03000001";
end if;
if first_state_sram_input_id = 5413 then
	sram_write <= x"82D05504";
end if;
if first_state_sram_input_id = 5414 then
	sram_write <= x"02A00002";
end if;
if first_state_sram_input_id = 5415 then
	sram_write <= x"82CA54C4";
end if;
if first_state_sram_input_id = 5416 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 5417 then
	sram_write <= x"00480000";
end if;
if first_state_sram_input_id = 5418 then
	sram_write <= x"002E0000";
end if;
if first_state_sram_input_id = 5419 then
	sram_write <= x"03DC0014";
end if;
if first_state_sram_input_id = 5420 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 5421 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 5422 then
	sram_write <= x"82003A54";
end if;
if first_state_sram_input_id = 5423 then
	sram_write <= x"07DC0014";
end if;
if first_state_sram_input_id = 5424 then
	sram_write <= x"82005500";
end if;
if first_state_sram_input_id = 5425 then
	sram_write <= x"C8880000";
end if;
if first_state_sram_input_id = 5426 then
	sram_write <= x"8E8054D4";
end if;
if first_state_sram_input_id = 5427 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 5428 then
	sram_write <= x"82005500";
end if;
if first_state_sram_input_id = 5429 then
	sram_write <= x"02A002AC";
end if;
if first_state_sram_input_id = 5430 then
	sram_write <= x"C8880004";
end if;
if first_state_sram_input_id = 5431 then
	sram_write <= x"48282000";
end if;
if first_state_sram_input_id = 5432 then
	sram_write <= x"C8880008";
end if;
if first_state_sram_input_id = 5433 then
	sram_write <= x"48484000";
end if;
if first_state_sram_input_id = 5434 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 5435 then
	sram_write <= x"C848000C";
end if;
if first_state_sram_input_id = 5436 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 5437 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 5438 then
	sram_write <= x"CC2A0000";
end if;
if first_state_sram_input_id = 5439 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 5440 then
	sram_write <= x"8200552C";
end if;
if first_state_sram_input_id = 5441 then
	sram_write <= x"C0AA0000";
end if;
if first_state_sram_input_id = 5442 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 5443 then
	sram_write <= x"00680000";
end if;
if first_state_sram_input_id = 5444 then
	sram_write <= x"004A0000";
end if;
if first_state_sram_input_id = 5445 then
	sram_write <= x"002E0000";
end if;
if first_state_sram_input_id = 5446 then
	sram_write <= x"03DC0014";
end if;
if first_state_sram_input_id = 5447 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 5448 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 5449 then
	sram_write <= x"8200389C";
end if;
if first_state_sram_input_id = 5450 then
	sram_write <= x"07DC0014";
end if;
if first_state_sram_input_id = 5451 then
	sram_write <= x"82205670";
end if;
if first_state_sram_input_id = 5452 then
	sram_write <= x"022002AC";
end if;
if first_state_sram_input_id = 5453 then
	sram_write <= x"C8220000";
end if;
if first_state_sram_input_id = 5454 then
	sram_write <= x"C8400070";
end if;
if first_state_sram_input_id = 5455 then
	sram_write <= x"8E245548";
end if;
if first_state_sram_input_id = 5456 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 5457 then
	sram_write <= x"8200566C";
end if;
if first_state_sram_input_id = 5458 then
	sram_write <= x"C03C0000";
end if;
if first_state_sram_input_id = 5459 then
	sram_write <= x"C0420004";
end if;
if first_state_sram_input_id = 5460 then
	sram_write <= x"0260FFFF";
end if;
if first_state_sram_input_id = 5461 then
	sram_write <= x"82465658";
end if;
if first_state_sram_input_id = 5462 then
	sram_write <= x"026001E0";
end if;
if first_state_sram_input_id = 5463 then
	sram_write <= x"22440220";
end if;
if first_state_sram_input_id = 5464 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 5465 then
	sram_write <= x"02800000";
end if;
if first_state_sram_input_id = 5466 then
	sram_write <= x"C47C000C";
end if;
if first_state_sram_input_id = 5467 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 5468 then
	sram_write <= x"00280000";
end if;
if first_state_sram_input_id = 5469 then
	sram_write <= x"03DC0018";
end if;
if first_state_sram_input_id = 5470 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 5471 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 5472 then
	sram_write <= x"82004E40";
end if;
if first_state_sram_input_id = 5473 then
	sram_write <= x"07DC0018";
end if;
if first_state_sram_input_id = 5474 then
	sram_write <= x"82205594";
end if;
if first_state_sram_input_id = 5475 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 5476 then
	sram_write <= x"82005654";
end if;
if first_state_sram_input_id = 5477 then
	sram_write <= x"C03C0000";
end if;
if first_state_sram_input_id = 5478 then
	sram_write <= x"C0420008";
end if;
if first_state_sram_input_id = 5479 then
	sram_write <= x"0260FFFF";
end if;
if first_state_sram_input_id = 5480 then
	sram_write <= x"82465650";
end if;
if first_state_sram_input_id = 5481 then
	sram_write <= x"22440220";
end if;
if first_state_sram_input_id = 5482 then
	sram_write <= x"C07C000C";
end if;
if first_state_sram_input_id = 5483 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 5484 then
	sram_write <= x"02800000";
end if;
if first_state_sram_input_id = 5485 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 5486 then
	sram_write <= x"00280000";
end if;
if first_state_sram_input_id = 5487 then
	sram_write <= x"03DC0018";
end if;
if first_state_sram_input_id = 5488 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 5489 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 5490 then
	sram_write <= x"82004E40";
end if;
if first_state_sram_input_id = 5491 then
	sram_write <= x"07DC0018";
end if;
if first_state_sram_input_id = 5492 then
	sram_write <= x"822055DC";
end if;
if first_state_sram_input_id = 5493 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 5494 then
	sram_write <= x"8200564C";
end if;
if first_state_sram_input_id = 5495 then
	sram_write <= x"C03C0000";
end if;
if first_state_sram_input_id = 5496 then
	sram_write <= x"C042000C";
end if;
if first_state_sram_input_id = 5497 then
	sram_write <= x"0260FFFF";
end if;
if first_state_sram_input_id = 5498 then
	sram_write <= x"82465648";
end if;
if first_state_sram_input_id = 5499 then
	sram_write <= x"22440220";
end if;
if first_state_sram_input_id = 5500 then
	sram_write <= x"C07C000C";
end if;
if first_state_sram_input_id = 5501 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 5502 then
	sram_write <= x"02600000";
end if;
if first_state_sram_input_id = 5503 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 5504 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 5505 then
	sram_write <= x"03DC0018";
end if;
if first_state_sram_input_id = 5506 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 5507 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 5508 then
	sram_write <= x"82004E40";
end if;
if first_state_sram_input_id = 5509 then
	sram_write <= x"07DC0018";
end if;
if first_state_sram_input_id = 5510 then
	sram_write <= x"82205624";
end if;
if first_state_sram_input_id = 5511 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 5512 then
	sram_write <= x"82005644";
end if;
if first_state_sram_input_id = 5513 then
	sram_write <= x"02200004";
end if;
if first_state_sram_input_id = 5514 then
	sram_write <= x"C05C0000";
end if;
if first_state_sram_input_id = 5515 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 5516 then
	sram_write <= x"03DC0018";
end if;
if first_state_sram_input_id = 5517 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 5518 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 5519 then
	sram_write <= x"82005284";
end if;
if first_state_sram_input_id = 5520 then
	sram_write <= x"07DC0018";
end if;
if first_state_sram_input_id = 5521 then
	sram_write <= x"8200564C";
end if;
if first_state_sram_input_id = 5522 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 5523 then
	sram_write <= x"82005654";
end if;
if first_state_sram_input_id = 5524 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 5525 then
	sram_write <= x"8200565C";
end if;
if first_state_sram_input_id = 5526 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 5527 then
	sram_write <= x"82205668";
end if;
if first_state_sram_input_id = 5528 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 5529 then
	sram_write <= x"8200566C";
end if;
if first_state_sram_input_id = 5530 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 5531 then
	sram_write <= x"82005674";
end if;
if first_state_sram_input_id = 5532 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 5533 then
	sram_write <= x"8200567C";
end if;
if first_state_sram_input_id = 5534 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 5535 then
	sram_write <= x"822057B0";
end if;
if first_state_sram_input_id = 5536 then
	sram_write <= x"C03C0000";
end if;
if first_state_sram_input_id = 5537 then
	sram_write <= x"C0420004";
end if;
if first_state_sram_input_id = 5538 then
	sram_write <= x"0260FFFF";
end if;
if first_state_sram_input_id = 5539 then
	sram_write <= x"82465790";
end if;
if first_state_sram_input_id = 5540 then
	sram_write <= x"026001E0";
end if;
if first_state_sram_input_id = 5541 then
	sram_write <= x"22440220";
end if;
if first_state_sram_input_id = 5542 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 5543 then
	sram_write <= x"02800000";
end if;
if first_state_sram_input_id = 5544 then
	sram_write <= x"C47C0010";
end if;
if first_state_sram_input_id = 5545 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 5546 then
	sram_write <= x"00280000";
end if;
if first_state_sram_input_id = 5547 then
	sram_write <= x"03DC001C";
end if;
if first_state_sram_input_id = 5548 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 5549 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 5550 then
	sram_write <= x"82004E40";
end if;
if first_state_sram_input_id = 5551 then
	sram_write <= x"07DC001C";
end if;
if first_state_sram_input_id = 5552 then
	sram_write <= x"822056CC";
end if;
if first_state_sram_input_id = 5553 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 5554 then
	sram_write <= x"8200578C";
end if;
if first_state_sram_input_id = 5555 then
	sram_write <= x"C03C0000";
end if;
if first_state_sram_input_id = 5556 then
	sram_write <= x"C0420008";
end if;
if first_state_sram_input_id = 5557 then
	sram_write <= x"0260FFFF";
end if;
if first_state_sram_input_id = 5558 then
	sram_write <= x"82465788";
end if;
if first_state_sram_input_id = 5559 then
	sram_write <= x"22440220";
end if;
if first_state_sram_input_id = 5560 then
	sram_write <= x"C07C0010";
end if;
if first_state_sram_input_id = 5561 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 5562 then
	sram_write <= x"02800000";
end if;
if first_state_sram_input_id = 5563 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 5564 then
	sram_write <= x"00280000";
end if;
if first_state_sram_input_id = 5565 then
	sram_write <= x"03DC001C";
end if;
if first_state_sram_input_id = 5566 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 5567 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 5568 then
	sram_write <= x"82004E40";
end if;
if first_state_sram_input_id = 5569 then
	sram_write <= x"07DC001C";
end if;
if first_state_sram_input_id = 5570 then
	sram_write <= x"82205714";
end if;
if first_state_sram_input_id = 5571 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 5572 then
	sram_write <= x"82005784";
end if;
if first_state_sram_input_id = 5573 then
	sram_write <= x"C03C0000";
end if;
if first_state_sram_input_id = 5574 then
	sram_write <= x"C042000C";
end if;
if first_state_sram_input_id = 5575 then
	sram_write <= x"0260FFFF";
end if;
if first_state_sram_input_id = 5576 then
	sram_write <= x"82465780";
end if;
if first_state_sram_input_id = 5577 then
	sram_write <= x"22440220";
end if;
if first_state_sram_input_id = 5578 then
	sram_write <= x"C07C0010";
end if;
if first_state_sram_input_id = 5579 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 5580 then
	sram_write <= x"02600000";
end if;
if first_state_sram_input_id = 5581 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 5582 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 5583 then
	sram_write <= x"03DC001C";
end if;
if first_state_sram_input_id = 5584 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 5585 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 5586 then
	sram_write <= x"82004E40";
end if;
if first_state_sram_input_id = 5587 then
	sram_write <= x"07DC001C";
end if;
if first_state_sram_input_id = 5588 then
	sram_write <= x"8220575C";
end if;
if first_state_sram_input_id = 5589 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 5590 then
	sram_write <= x"8200577C";
end if;
if first_state_sram_input_id = 5591 then
	sram_write <= x"02200004";
end if;
if first_state_sram_input_id = 5592 then
	sram_write <= x"C05C0000";
end if;
if first_state_sram_input_id = 5593 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 5594 then
	sram_write <= x"03DC001C";
end if;
if first_state_sram_input_id = 5595 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 5596 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 5597 then
	sram_write <= x"82005284";
end if;
if first_state_sram_input_id = 5598 then
	sram_write <= x"07DC001C";
end if;
if first_state_sram_input_id = 5599 then
	sram_write <= x"82005784";
end if;
if first_state_sram_input_id = 5600 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 5601 then
	sram_write <= x"8200578C";
end if;
if first_state_sram_input_id = 5602 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 5603 then
	sram_write <= x"82005794";
end if;
if first_state_sram_input_id = 5604 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 5605 then
	sram_write <= x"822057A0";
end if;
if first_state_sram_input_id = 5606 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 5607 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 5608 then
	sram_write <= x"C03C0008";
end if;
if first_state_sram_input_id = 5609 then
	sram_write <= x"02220001";
end if;
if first_state_sram_input_id = 5610 then
	sram_write <= x"C05C0004";
end if;
if first_state_sram_input_id = 5611 then
	sram_write <= x"82005414";
end if;
if first_state_sram_input_id = 5612 then
	sram_write <= x"C03C0008";
end if;
if first_state_sram_input_id = 5613 then
	sram_write <= x"02220001";
end if;
if first_state_sram_input_id = 5614 then
	sram_write <= x"C05C0004";
end if;
if first_state_sram_input_id = 5615 then
	sram_write <= x"82005414";
end if;
if first_state_sram_input_id = 5616 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 5617 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 5618 then
	sram_write <= x"22820220";
end if;
if first_state_sram_input_id = 5619 then
	sram_write <= x"D0848000";
end if;
if first_state_sram_input_id = 5620 then
	sram_write <= x"02A0FFFF";
end if;
if first_state_sram_input_id = 5621 then
	sram_write <= x"828A5CD8";
end if;
if first_state_sram_input_id = 5622 then
	sram_write <= x"02A0030C";
end if;
if first_state_sram_input_id = 5623 then
	sram_write <= x"02C000C8";
end if;
if first_state_sram_input_id = 5624 then
	sram_write <= x"22E80220";
end if;
if first_state_sram_input_id = 5625 then
	sram_write <= x"D0ECE000";
end if;
if first_state_sram_input_id = 5626 then
	sram_write <= x"C82A0000";
end if;
if first_state_sram_input_id = 5627 then
	sram_write <= x"C10E0014";
end if;
if first_state_sram_input_id = 5628 then
	sram_write <= x"C8500000";
end if;
if first_state_sram_input_id = 5629 then
	sram_write <= x"44224000";
end if;
if first_state_sram_input_id = 5630 then
	sram_write <= x"C84A0004";
end if;
if first_state_sram_input_id = 5631 then
	sram_write <= x"C10E0014";
end if;
if first_state_sram_input_id = 5632 then
	sram_write <= x"C8700004";
end if;
if first_state_sram_input_id = 5633 then
	sram_write <= x"44446000";
end if;
if first_state_sram_input_id = 5634 then
	sram_write <= x"C86A0008";
end if;
if first_state_sram_input_id = 5635 then
	sram_write <= x"C10E0014";
end if;
if first_state_sram_input_id = 5636 then
	sram_write <= x"C8900008";
end if;
if first_state_sram_input_id = 5637 then
	sram_write <= x"44668000";
end if;
if first_state_sram_input_id = 5638 then
	sram_write <= x"C10E0004";
end if;
if first_state_sram_input_id = 5639 then
	sram_write <= x"03200001";
end if;
if first_state_sram_input_id = 5640 then
	sram_write <= x"C4BC0000";
end if;
if first_state_sram_input_id = 5641 then
	sram_write <= x"C47C0004";
end if;
if first_state_sram_input_id = 5642 then
	sram_write <= x"C45C0008";
end if;
if first_state_sram_input_id = 5643 then
	sram_write <= x"C43C000C";
end if;
if first_state_sram_input_id = 5644 then
	sram_write <= x"C4DC0010";
end if;
if first_state_sram_input_id = 5645 then
	sram_write <= x"C49C0014";
end if;
if first_state_sram_input_id = 5646 then
	sram_write <= x"8312588C";
end if;
if first_state_sram_input_id = 5647 then
	sram_write <= x"03200002";
end if;
if first_state_sram_input_id = 5648 then
	sram_write <= x"83125868";
end if;
if first_state_sram_input_id = 5649 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 5650 then
	sram_write <= x"00460000";
end if;
if first_state_sram_input_id = 5651 then
	sram_write <= x"002E0000";
end if;
if first_state_sram_input_id = 5652 then
	sram_write <= x"03DC0020";
end if;
if first_state_sram_input_id = 5653 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 5654 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 5655 then
	sram_write <= x"820034A0";
end if;
if first_state_sram_input_id = 5656 then
	sram_write <= x"07DC0020";
end if;
if first_state_sram_input_id = 5657 then
	sram_write <= x"82005888";
end if;
if first_state_sram_input_id = 5658 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 5659 then
	sram_write <= x"00460000";
end if;
if first_state_sram_input_id = 5660 then
	sram_write <= x"002E0000";
end if;
if first_state_sram_input_id = 5661 then
	sram_write <= x"03DC0020";
end if;
if first_state_sram_input_id = 5662 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 5663 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 5664 then
	sram_write <= x"820032A4";
end if;
if first_state_sram_input_id = 5665 then
	sram_write <= x"07DC0020";
end if;
if first_state_sram_input_id = 5666 then
	sram_write <= x"8200596C";
end if;
if first_state_sram_input_id = 5667 then
	sram_write <= x"03000000";
end if;
if first_state_sram_input_id = 5668 then
	sram_write <= x"03200001";
end if;
if first_state_sram_input_id = 5669 then
	sram_write <= x"03400002";
end if;
if first_state_sram_input_id = 5670 then
	sram_write <= x"CC3C0018";
end if;
if first_state_sram_input_id = 5671 then
	sram_write <= x"CC7C0020";
end if;
if first_state_sram_input_id = 5672 then
	sram_write <= x"CC5C0028";
end if;
if first_state_sram_input_id = 5673 then
	sram_write <= x"C4FC0030";
end if;
if first_state_sram_input_id = 5674 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 5675 then
	sram_write <= x"00B40000";
end if;
if first_state_sram_input_id = 5676 then
	sram_write <= x"00920000";
end if;
if first_state_sram_input_id = 5677 then
	sram_write <= x"00460000";
end if;
if first_state_sram_input_id = 5678 then
	sram_write <= x"002E0000";
end if;
if first_state_sram_input_id = 5679 then
	sram_write <= x"00700000";
end if;
if first_state_sram_input_id = 5680 then
	sram_write <= x"03DC003C";
end if;
if first_state_sram_input_id = 5681 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 5682 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 5683 then
	sram_write <= x"8200317C";
end if;
if first_state_sram_input_id = 5684 then
	sram_write <= x"07DC003C";
end if;
if first_state_sram_input_id = 5685 then
	sram_write <= x"822058E0";
end if;
if first_state_sram_input_id = 5686 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 5687 then
	sram_write <= x"8200596C";
end if;
if first_state_sram_input_id = 5688 then
	sram_write <= x"02600001";
end if;
if first_state_sram_input_id = 5689 then
	sram_write <= x"02800002";
end if;
if first_state_sram_input_id = 5690 then
	sram_write <= x"02A00000";
end if;
if first_state_sram_input_id = 5691 then
	sram_write <= x"C83C0028";
end if;
if first_state_sram_input_id = 5692 then
	sram_write <= x"C85C0020";
end if;
if first_state_sram_input_id = 5693 then
	sram_write <= x"C87C0018";
end if;
if first_state_sram_input_id = 5694 then
	sram_write <= x"C03C0030";
end if;
if first_state_sram_input_id = 5695 then
	sram_write <= x"C05C0004";
end if;
if first_state_sram_input_id = 5696 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 5697 then
	sram_write <= x"03DC003C";
end if;
if first_state_sram_input_id = 5698 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 5699 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 5700 then
	sram_write <= x"8200317C";
end if;
if first_state_sram_input_id = 5701 then
	sram_write <= x"07DC003C";
end if;
if first_state_sram_input_id = 5702 then
	sram_write <= x"82205924";
end if;
if first_state_sram_input_id = 5703 then
	sram_write <= x"02200002";
end if;
if first_state_sram_input_id = 5704 then
	sram_write <= x"8200596C";
end if;
if first_state_sram_input_id = 5705 then
	sram_write <= x"02600002";
end if;
if first_state_sram_input_id = 5706 then
	sram_write <= x"02800000";
end if;
if first_state_sram_input_id = 5707 then
	sram_write <= x"02A00001";
end if;
if first_state_sram_input_id = 5708 then
	sram_write <= x"C83C0020";
end if;
if first_state_sram_input_id = 5709 then
	sram_write <= x"C85C0018";
end if;
if first_state_sram_input_id = 5710 then
	sram_write <= x"C87C0028";
end if;
if first_state_sram_input_id = 5711 then
	sram_write <= x"C03C0030";
end if;
if first_state_sram_input_id = 5712 then
	sram_write <= x"C05C0004";
end if;
if first_state_sram_input_id = 5713 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 5714 then
	sram_write <= x"03DC003C";
end if;
if first_state_sram_input_id = 5715 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 5716 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 5717 then
	sram_write <= x"8200317C";
end if;
if first_state_sram_input_id = 5718 then
	sram_write <= x"07DC003C";
end if;
if first_state_sram_input_id = 5719 then
	sram_write <= x"82205968";
end if;
if first_state_sram_input_id = 5720 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 5721 then
	sram_write <= x"8200596C";
end if;
if first_state_sram_input_id = 5722 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 5723 then
	sram_write <= x"82205CA8";
end if;
if first_state_sram_input_id = 5724 then
	sram_write <= x"024002AC";
end if;
if first_state_sram_input_id = 5725 then
	sram_write <= x"C8240000";
end if;
if first_state_sram_input_id = 5726 then
	sram_write <= x"8E025980";
end if;
if first_state_sram_input_id = 5727 then
	sram_write <= x"82005C94";
end if;
if first_state_sram_input_id = 5728 then
	sram_write <= x"024002B4";
end if;
if first_state_sram_input_id = 5729 then
	sram_write <= x"C8440000";
end if;
if first_state_sram_input_id = 5730 then
	sram_write <= x"8E245990";
end if;
if first_state_sram_input_id = 5731 then
	sram_write <= x"82005C94";
end if;
if first_state_sram_input_id = 5732 then
	sram_write <= x"C8400074";
end if;
if first_state_sram_input_id = 5733 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 5734 then
	sram_write <= x"C07C0004";
end if;
if first_state_sram_input_id = 5735 then
	sram_write <= x"C8460000";
end if;
if first_state_sram_input_id = 5736 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 5737 then
	sram_write <= x"C09C0000";
end if;
if first_state_sram_input_id = 5738 then
	sram_write <= x"C8680000";
end if;
if first_state_sram_input_id = 5739 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 5740 then
	sram_write <= x"C8660004";
end if;
if first_state_sram_input_id = 5741 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 5742 then
	sram_write <= x"C8880004";
end if;
if first_state_sram_input_id = 5743 then
	sram_write <= x"40668000";
end if;
if first_state_sram_input_id = 5744 then
	sram_write <= x"C8860008";
end if;
if first_state_sram_input_id = 5745 then
	sram_write <= x"48882000";
end if;
if first_state_sram_input_id = 5746 then
	sram_write <= x"C8A80008";
end if;
if first_state_sram_input_id = 5747 then
	sram_write <= x"4088A000";
end if;
if first_state_sram_input_id = 5748 then
	sram_write <= x"C09C0008";
end if;
if first_state_sram_input_id = 5749 then
	sram_write <= x"C0A80000";
end if;
if first_state_sram_input_id = 5750 then
	sram_write <= x"02C0FFFF";
end if;
if first_state_sram_input_id = 5751 then
	sram_write <= x"C43C0034";
end if;
if first_state_sram_input_id = 5752 then
	sram_write <= x"CC9C0038";
end if;
if first_state_sram_input_id = 5753 then
	sram_write <= x"CC7C0040";
end if;
if first_state_sram_input_id = 5754 then
	sram_write <= x"CC5C0048";
end if;
if first_state_sram_input_id = 5755 then
	sram_write <= x"C45C0050";
end if;
if first_state_sram_input_id = 5756 then
	sram_write <= x"CC3C0058";
end if;
if first_state_sram_input_id = 5757 then
	sram_write <= x"82AC5C48";
end if;
if first_state_sram_input_id = 5758 then
	sram_write <= x"22AA0220";
end if;
if first_state_sram_input_id = 5759 then
	sram_write <= x"C0DC0010";
end if;
if first_state_sram_input_id = 5760 then
	sram_write <= x"D0ACA000";
end if;
if first_state_sram_input_id = 5761 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 5762 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 5763 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 5764 then
	sram_write <= x"40406000";
end if;
if first_state_sram_input_id = 5765 then
	sram_write <= x"40608000";
end if;
if first_state_sram_input_id = 5766 then
	sram_write <= x"03DC0068";
end if;
if first_state_sram_input_id = 5767 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 5768 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 5769 then
	sram_write <= x"82004860";
end if;
if first_state_sram_input_id = 5770 then
	sram_write <= x"07DC0068";
end if;
if first_state_sram_input_id = 5771 then
	sram_write <= x"82205A38";
end if;
if first_state_sram_input_id = 5772 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 5773 then
	sram_write <= x"82005C44";
end if;
if first_state_sram_input_id = 5774 then
	sram_write <= x"C05C0008";
end if;
if first_state_sram_input_id = 5775 then
	sram_write <= x"C0240004";
end if;
if first_state_sram_input_id = 5776 then
	sram_write <= x"0260FFFF";
end if;
if first_state_sram_input_id = 5777 then
	sram_write <= x"82265C40";
end if;
if first_state_sram_input_id = 5778 then
	sram_write <= x"22220220";
end if;
if first_state_sram_input_id = 5779 then
	sram_write <= x"C07C0010";
end if;
if first_state_sram_input_id = 5780 then
	sram_write <= x"D0262000";
end if;
if first_state_sram_input_id = 5781 then
	sram_write <= x"C0820014";
end if;
if first_state_sram_input_id = 5782 then
	sram_write <= x"C8280000";
end if;
if first_state_sram_input_id = 5783 then
	sram_write <= x"C85C0048";
end if;
if first_state_sram_input_id = 5784 then
	sram_write <= x"44242000";
end if;
if first_state_sram_input_id = 5785 then
	sram_write <= x"C0820014";
end if;
if first_state_sram_input_id = 5786 then
	sram_write <= x"C8680004";
end if;
if first_state_sram_input_id = 5787 then
	sram_write <= x"C89C0040";
end if;
if first_state_sram_input_id = 5788 then
	sram_write <= x"44686000";
end if;
if first_state_sram_input_id = 5789 then
	sram_write <= x"C0820014";
end if;
if first_state_sram_input_id = 5790 then
	sram_write <= x"C8A80008";
end if;
if first_state_sram_input_id = 5791 then
	sram_write <= x"C8DC0038";
end if;
if first_state_sram_input_id = 5792 then
	sram_write <= x"44ACA000";
end if;
if first_state_sram_input_id = 5793 then
	sram_write <= x"C0820004";
end if;
if first_state_sram_input_id = 5794 then
	sram_write <= x"02A00001";
end if;
if first_state_sram_input_id = 5795 then
	sram_write <= x"828A5B24";
end if;
if first_state_sram_input_id = 5796 then
	sram_write <= x"02A00002";
end if;
if first_state_sram_input_id = 5797 then
	sram_write <= x"828A5ABC";
end if;
if first_state_sram_input_id = 5798 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 5799 then
	sram_write <= x"40406000";
end if;
if first_state_sram_input_id = 5800 then
	sram_write <= x"4060A000";
end if;
if first_state_sram_input_id = 5801 then
	sram_write <= x"03DC0068";
end if;
if first_state_sram_input_id = 5802 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 5803 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 5804 then
	sram_write <= x"82004780";
end if;
if first_state_sram_input_id = 5805 then
	sram_write <= x"07DC0068";
end if;
if first_state_sram_input_id = 5806 then
	sram_write <= x"82005B20";
end if;
if first_state_sram_input_id = 5807 then
	sram_write <= x"C0820010";
end if;
if first_state_sram_input_id = 5808 then
	sram_write <= x"C8E80000";
end if;
if first_state_sram_input_id = 5809 then
	sram_write <= x"482E2000";
end if;
if first_state_sram_input_id = 5810 then
	sram_write <= x"C8E80004";
end if;
if first_state_sram_input_id = 5811 then
	sram_write <= x"486E6000";
end if;
if first_state_sram_input_id = 5812 then
	sram_write <= x"40226000";
end if;
if first_state_sram_input_id = 5813 then
	sram_write <= x"C8680008";
end if;
if first_state_sram_input_id = 5814 then
	sram_write <= x"4866A000";
end if;
if first_state_sram_input_id = 5815 then
	sram_write <= x"40226000";
end if;
if first_state_sram_input_id = 5816 then
	sram_write <= x"C0220018";
end if;
if first_state_sram_input_id = 5817 then
	sram_write <= x"8E205AF0";
end if;
if first_state_sram_input_id = 5818 then
	sram_write <= x"02800000";
end if;
if first_state_sram_input_id = 5819 then
	sram_write <= x"82005AF4";
end if;
if first_state_sram_input_id = 5820 then
	sram_write <= x"02800001";
end if;
if first_state_sram_input_id = 5821 then
	sram_write <= x"82205B0C";
end if;
if first_state_sram_input_id = 5822 then
	sram_write <= x"8E205B04";
end if;
if first_state_sram_input_id = 5823 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 5824 then
	sram_write <= x"82005B08";
end if;
if first_state_sram_input_id = 5825 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 5826 then
	sram_write <= x"82005B10";
end if;
if first_state_sram_input_id = 5827 then
	sram_write <= x"00280000";
end if;
if first_state_sram_input_id = 5828 then
	sram_write <= x"82205B1C";
end if;
if first_state_sram_input_id = 5829 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 5830 then
	sram_write <= x"82005B20";
end if;
if first_state_sram_input_id = 5831 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 5832 then
	sram_write <= x"82005BB0";
end if;
if first_state_sram_input_id = 5833 then
	sram_write <= x"8E205B2C";
end if;
if first_state_sram_input_id = 5834 then
	sram_write <= x"82005B30";
end if;
if first_state_sram_input_id = 5835 then
	sram_write <= x"44202000";
end if;
if first_state_sram_input_id = 5836 then
	sram_write <= x"C0820010";
end if;
if first_state_sram_input_id = 5837 then
	sram_write <= x"C8E80000";
end if;
if first_state_sram_input_id = 5838 then
	sram_write <= x"8E2E5B44";
end if;
if first_state_sram_input_id = 5839 then
	sram_write <= x"02800000";
end if;
if first_state_sram_input_id = 5840 then
	sram_write <= x"82005B90";
end if;
if first_state_sram_input_id = 5841 then
	sram_write <= x"8E605B50";
end if;
if first_state_sram_input_id = 5842 then
	sram_write <= x"40206000";
end if;
if first_state_sram_input_id = 5843 then
	sram_write <= x"82005B54";
end if;
if first_state_sram_input_id = 5844 then
	sram_write <= x"44206000";
end if;
if first_state_sram_input_id = 5845 then
	sram_write <= x"C0820010";
end if;
if first_state_sram_input_id = 5846 then
	sram_write <= x"C8680004";
end if;
if first_state_sram_input_id = 5847 then
	sram_write <= x"8E265B68";
end if;
if first_state_sram_input_id = 5848 then
	sram_write <= x"02800000";
end if;
if first_state_sram_input_id = 5849 then
	sram_write <= x"82005B90";
end if;
if first_state_sram_input_id = 5850 then
	sram_write <= x"8EA05B74";
end if;
if first_state_sram_input_id = 5851 then
	sram_write <= x"4020A000";
end if;
if first_state_sram_input_id = 5852 then
	sram_write <= x"82005B78";
end if;
if first_state_sram_input_id = 5853 then
	sram_write <= x"4420A000";
end if;
if first_state_sram_input_id = 5854 then
	sram_write <= x"C0820010";
end if;
if first_state_sram_input_id = 5855 then
	sram_write <= x"C8680008";
end if;
if first_state_sram_input_id = 5856 then
	sram_write <= x"8E265B8C";
end if;
if first_state_sram_input_id = 5857 then
	sram_write <= x"02800000";
end if;
if first_state_sram_input_id = 5858 then
	sram_write <= x"82005B90";
end if;
if first_state_sram_input_id = 5859 then
	sram_write <= x"02800001";
end if;
if first_state_sram_input_id = 5860 then
	sram_write <= x"82805B9C";
end if;
if first_state_sram_input_id = 5861 then
	sram_write <= x"C0220018";
end if;
if first_state_sram_input_id = 5862 then
	sram_write <= x"82005BB0";
end if;
if first_state_sram_input_id = 5863 then
	sram_write <= x"C0220018";
end if;
if first_state_sram_input_id = 5864 then
	sram_write <= x"82205BAC";
end if;
if first_state_sram_input_id = 5865 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 5866 then
	sram_write <= x"82005BB0";
end if;
if first_state_sram_input_id = 5867 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 5868 then
	sram_write <= x"82205BBC";
end if;
if first_state_sram_input_id = 5869 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 5870 then
	sram_write <= x"82005C3C";
end if;
if first_state_sram_input_id = 5871 then
	sram_write <= x"C05C0008";
end if;
if first_state_sram_input_id = 5872 then
	sram_write <= x"C0240008";
end if;
if first_state_sram_input_id = 5873 then
	sram_write <= x"0260FFFF";
end if;
if first_state_sram_input_id = 5874 then
	sram_write <= x"82265C38";
end if;
if first_state_sram_input_id = 5875 then
	sram_write <= x"22220220";
end if;
if first_state_sram_input_id = 5876 then
	sram_write <= x"C07C0010";
end if;
if first_state_sram_input_id = 5877 then
	sram_write <= x"D0262000";
end if;
if first_state_sram_input_id = 5878 then
	sram_write <= x"C83C0048";
end if;
if first_state_sram_input_id = 5879 then
	sram_write <= x"C85C0040";
end if;
if first_state_sram_input_id = 5880 then
	sram_write <= x"C87C0038";
end if;
if first_state_sram_input_id = 5881 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 5882 then
	sram_write <= x"03DC0068";
end if;
if first_state_sram_input_id = 5883 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 5884 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 5885 then
	sram_write <= x"82004860";
end if;
if first_state_sram_input_id = 5886 then
	sram_write <= x"07DC0068";
end if;
if first_state_sram_input_id = 5887 then
	sram_write <= x"82205C08";
end if;
if first_state_sram_input_id = 5888 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 5889 then
	sram_write <= x"82005C34";
end if;
if first_state_sram_input_id = 5890 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 5891 then
	sram_write <= x"C83C0048";
end if;
if first_state_sram_input_id = 5892 then
	sram_write <= x"C85C0040";
end if;
if first_state_sram_input_id = 5893 then
	sram_write <= x"C87C0038";
end if;
if first_state_sram_input_id = 5894 then
	sram_write <= x"C05C0008";
end if;
if first_state_sram_input_id = 5895 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 5896 then
	sram_write <= x"03DC0068";
end if;
if first_state_sram_input_id = 5897 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 5898 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 5899 then
	sram_write <= x"82004A0C";
end if;
if first_state_sram_input_id = 5900 then
	sram_write <= x"07DC0068";
end if;
if first_state_sram_input_id = 5901 then
	sram_write <= x"82005C3C";
end if;
if first_state_sram_input_id = 5902 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 5903 then
	sram_write <= x"82005C44";
end if;
if first_state_sram_input_id = 5904 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 5905 then
	sram_write <= x"82005C4C";
end if;
if first_state_sram_input_id = 5906 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 5907 then
	sram_write <= x"82205C94";
end if;
if first_state_sram_input_id = 5908 then
	sram_write <= x"C03C0050";
end if;
if first_state_sram_input_id = 5909 then
	sram_write <= x"C83C0058";
end if;
if first_state_sram_input_id = 5910 then
	sram_write <= x"CC220000";
end if;
if first_state_sram_input_id = 5911 then
	sram_write <= x"022002B8";
end if;
if first_state_sram_input_id = 5912 then
	sram_write <= x"C83C0048";
end if;
if first_state_sram_input_id = 5913 then
	sram_write <= x"CC220000";
end if;
if first_state_sram_input_id = 5914 then
	sram_write <= x"C83C0040";
end if;
if first_state_sram_input_id = 5915 then
	sram_write <= x"CC220004";
end if;
if first_state_sram_input_id = 5916 then
	sram_write <= x"C83C0038";
end if;
if first_state_sram_input_id = 5917 then
	sram_write <= x"CC220008";
end if;
if first_state_sram_input_id = 5918 then
	sram_write <= x"022002C4";
end if;
if first_state_sram_input_id = 5919 then
	sram_write <= x"C05C0014";
end if;
if first_state_sram_input_id = 5920 then
	sram_write <= x"C4420000";
end if;
if first_state_sram_input_id = 5921 then
	sram_write <= x"022002B0";
end if;
if first_state_sram_input_id = 5922 then
	sram_write <= x"C05C0034";
end if;
if first_state_sram_input_id = 5923 then
	sram_write <= x"C4420000";
end if;
if first_state_sram_input_id = 5924 then
	sram_write <= x"82005C94";
end if;
if first_state_sram_input_id = 5925 then
	sram_write <= x"C03C000C";
end if;
if first_state_sram_input_id = 5926 then
	sram_write <= x"02220001";
end if;
if first_state_sram_input_id = 5927 then
	sram_write <= x"C05C0008";
end if;
if first_state_sram_input_id = 5928 then
	sram_write <= x"C07C0004";
end if;
if first_state_sram_input_id = 5929 then
	sram_write <= x"820057C8";
end if;
if first_state_sram_input_id = 5930 then
	sram_write <= x"C03C0014";
end if;
if first_state_sram_input_id = 5931 then
	sram_write <= x"22220220";
end if;
if first_state_sram_input_id = 5932 then
	sram_write <= x"C05C0010";
end if;
if first_state_sram_input_id = 5933 then
	sram_write <= x"D0242000";
end if;
if first_state_sram_input_id = 5934 then
	sram_write <= x"C0220018";
end if;
if first_state_sram_input_id = 5935 then
	sram_write <= x"82205CD4";
end if;
if first_state_sram_input_id = 5936 then
	sram_write <= x"C03C000C";
end if;
if first_state_sram_input_id = 5937 then
	sram_write <= x"02220001";
end if;
if first_state_sram_input_id = 5938 then
	sram_write <= x"C05C0008";
end if;
if first_state_sram_input_id = 5939 then
	sram_write <= x"C07C0004";
end if;
if first_state_sram_input_id = 5940 then
	sram_write <= x"820057C8";
end if;
if first_state_sram_input_id = 5941 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 5942 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 5943 then
	sram_write <= x"22820220";
end if;
if first_state_sram_input_id = 5944 then
	sram_write <= x"D0848000";
end if;
if first_state_sram_input_id = 5945 then
	sram_write <= x"02A0FFFF";
end if;
if first_state_sram_input_id = 5946 then
	sram_write <= x"828A5E48";
end if;
if first_state_sram_input_id = 5947 then
	sram_write <= x"02A001E0";
end if;
if first_state_sram_input_id = 5948 then
	sram_write <= x"22880220";
end if;
if first_state_sram_input_id = 5949 then
	sram_write <= x"D08A8000";
end if;
if first_state_sram_input_id = 5950 then
	sram_write <= x"02C00000";
end if;
if first_state_sram_input_id = 5951 then
	sram_write <= x"C47C0000";
end if;
if first_state_sram_input_id = 5952 then
	sram_write <= x"C4BC0004";
end if;
if first_state_sram_input_id = 5953 then
	sram_write <= x"C45C0008";
end if;
if first_state_sram_input_id = 5954 then
	sram_write <= x"C43C000C";
end if;
if first_state_sram_input_id = 5955 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 5956 then
	sram_write <= x"00480000";
end if;
if first_state_sram_input_id = 5957 then
	sram_write <= x"002C0000";
end if;
if first_state_sram_input_id = 5958 then
	sram_write <= x"03DC0018";
end if;
if first_state_sram_input_id = 5959 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 5960 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 5961 then
	sram_write <= x"820057C8";
end if;
if first_state_sram_input_id = 5962 then
	sram_write <= x"07DC0018";
end if;
if first_state_sram_input_id = 5963 then
	sram_write <= x"C03C000C";
end if;
if first_state_sram_input_id = 5964 then
	sram_write <= x"02220001";
end if;
if first_state_sram_input_id = 5965 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 5966 then
	sram_write <= x"C07C0008";
end if;
if first_state_sram_input_id = 5967 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 5968 then
	sram_write <= x"0280FFFF";
end if;
if first_state_sram_input_id = 5969 then
	sram_write <= x"82485E44";
end if;
if first_state_sram_input_id = 5970 then
	sram_write <= x"22440220";
end if;
if first_state_sram_input_id = 5971 then
	sram_write <= x"C09C0004";
end if;
if first_state_sram_input_id = 5972 then
	sram_write <= x"D0484000";
end if;
if first_state_sram_input_id = 5973 then
	sram_write <= x"02A00000";
end if;
if first_state_sram_input_id = 5974 then
	sram_write <= x"C0DC0000";
end if;
if first_state_sram_input_id = 5975 then
	sram_write <= x"C43C0010";
end if;
if first_state_sram_input_id = 5976 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 5977 then
	sram_write <= x"006C0000";
end if;
if first_state_sram_input_id = 5978 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 5979 then
	sram_write <= x"03DC001C";
end if;
if first_state_sram_input_id = 5980 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 5981 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 5982 then
	sram_write <= x"820057C8";
end if;
if first_state_sram_input_id = 5983 then
	sram_write <= x"07DC001C";
end if;
if first_state_sram_input_id = 5984 then
	sram_write <= x"C03C0010";
end if;
if first_state_sram_input_id = 5985 then
	sram_write <= x"02220001";
end if;
if first_state_sram_input_id = 5986 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 5987 then
	sram_write <= x"C07C0008";
end if;
if first_state_sram_input_id = 5988 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 5989 then
	sram_write <= x"0280FFFF";
end if;
if first_state_sram_input_id = 5990 then
	sram_write <= x"82485E40";
end if;
if first_state_sram_input_id = 5991 then
	sram_write <= x"22440220";
end if;
if first_state_sram_input_id = 5992 then
	sram_write <= x"C09C0004";
end if;
if first_state_sram_input_id = 5993 then
	sram_write <= x"D0484000";
end if;
if first_state_sram_input_id = 5994 then
	sram_write <= x"02A00000";
end if;
if first_state_sram_input_id = 5995 then
	sram_write <= x"C0DC0000";
end if;
if first_state_sram_input_id = 5996 then
	sram_write <= x"C43C0014";
end if;
if first_state_sram_input_id = 5997 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 5998 then
	sram_write <= x"006C0000";
end if;
if first_state_sram_input_id = 5999 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 6000 then
	sram_write <= x"03DC0020";
end if;
if first_state_sram_input_id = 6001 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 6002 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 6003 then
	sram_write <= x"820057C8";
end if;
if first_state_sram_input_id = 6004 then
	sram_write <= x"07DC0020";
end if;
if first_state_sram_input_id = 6005 then
	sram_write <= x"C03C0014";
end if;
if first_state_sram_input_id = 6006 then
	sram_write <= x"02220001";
end if;
if first_state_sram_input_id = 6007 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 6008 then
	sram_write <= x"C07C0008";
end if;
if first_state_sram_input_id = 6009 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 6010 then
	sram_write <= x"0280FFFF";
end if;
if first_state_sram_input_id = 6011 then
	sram_write <= x"82485E3C";
end if;
if first_state_sram_input_id = 6012 then
	sram_write <= x"22440220";
end if;
if first_state_sram_input_id = 6013 then
	sram_write <= x"C09C0004";
end if;
if first_state_sram_input_id = 6014 then
	sram_write <= x"D0484000";
end if;
if first_state_sram_input_id = 6015 then
	sram_write <= x"02800000";
end if;
if first_state_sram_input_id = 6016 then
	sram_write <= x"C0BC0000";
end if;
if first_state_sram_input_id = 6017 then
	sram_write <= x"C43C0018";
end if;
if first_state_sram_input_id = 6018 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 6019 then
	sram_write <= x"006A0000";
end if;
if first_state_sram_input_id = 6020 then
	sram_write <= x"00280000";
end if;
if first_state_sram_input_id = 6021 then
	sram_write <= x"03DC0024";
end if;
if first_state_sram_input_id = 6022 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 6023 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 6024 then
	sram_write <= x"820057C8";
end if;
if first_state_sram_input_id = 6025 then
	sram_write <= x"07DC0024";
end if;
if first_state_sram_input_id = 6026 then
	sram_write <= x"C03C0018";
end if;
if first_state_sram_input_id = 6027 then
	sram_write <= x"02220001";
end if;
if first_state_sram_input_id = 6028 then
	sram_write <= x"C05C0008";
end if;
if first_state_sram_input_id = 6029 then
	sram_write <= x"C07C0000";
end if;
if first_state_sram_input_id = 6030 then
	sram_write <= x"82005CDC";
end if;
if first_state_sram_input_id = 6031 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 6032 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 6033 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 6034 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 6035 then
	sram_write <= x"22820220";
end if;
if first_state_sram_input_id = 6036 then
	sram_write <= x"D0848000";
end if;
if first_state_sram_input_id = 6037 then
	sram_write <= x"C0A80000";
end if;
if first_state_sram_input_id = 6038 then
	sram_write <= x"02C0FFFF";
end if;
if first_state_sram_input_id = 6039 then
	sram_write <= x"82AC6420";
end if;
if first_state_sram_input_id = 6040 then
	sram_write <= x"02C00063";
end if;
if first_state_sram_input_id = 6041 then
	sram_write <= x"C47C0000";
end if;
if first_state_sram_input_id = 6042 then
	sram_write <= x"C45C0004";
end if;
if first_state_sram_input_id = 6043 then
	sram_write <= x"C43C0008";
end if;
if first_state_sram_input_id = 6044 then
	sram_write <= x"82AC6118";
end if;
if first_state_sram_input_id = 6045 then
	sram_write <= x"02C0030C";
end if;
if first_state_sram_input_id = 6046 then
	sram_write <= x"02E000C8";
end if;
if first_state_sram_input_id = 6047 then
	sram_write <= x"22AA0220";
end if;
if first_state_sram_input_id = 6048 then
	sram_write <= x"D0AEA000";
end if;
if first_state_sram_input_id = 6049 then
	sram_write <= x"C82C0000";
end if;
if first_state_sram_input_id = 6050 then
	sram_write <= x"C0EA0014";
end if;
if first_state_sram_input_id = 6051 then
	sram_write <= x"C84E0000";
end if;
if first_state_sram_input_id = 6052 then
	sram_write <= x"44224000";
end if;
if first_state_sram_input_id = 6053 then
	sram_write <= x"C84C0004";
end if;
if first_state_sram_input_id = 6054 then
	sram_write <= x"C0EA0014";
end if;
if first_state_sram_input_id = 6055 then
	sram_write <= x"C86E0004";
end if;
if first_state_sram_input_id = 6056 then
	sram_write <= x"44446000";
end if;
if first_state_sram_input_id = 6057 then
	sram_write <= x"C86C0008";
end if;
if first_state_sram_input_id = 6058 then
	sram_write <= x"C0CA0014";
end if;
if first_state_sram_input_id = 6059 then
	sram_write <= x"C88C0008";
end if;
if first_state_sram_input_id = 6060 then
	sram_write <= x"44668000";
end if;
if first_state_sram_input_id = 6061 then
	sram_write <= x"C0CA0004";
end if;
if first_state_sram_input_id = 6062 then
	sram_write <= x"02E00001";
end if;
if first_state_sram_input_id = 6063 then
	sram_write <= x"C49C000C";
end if;
if first_state_sram_input_id = 6064 then
	sram_write <= x"82CE5F14";
end if;
if first_state_sram_input_id = 6065 then
	sram_write <= x"02E00002";
end if;
if first_state_sram_input_id = 6066 then
	sram_write <= x"82CE5EF0";
end if;
if first_state_sram_input_id = 6067 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 6068 then
	sram_write <= x"00460000";
end if;
if first_state_sram_input_id = 6069 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 6070 then
	sram_write <= x"03DC0018";
end if;
if first_state_sram_input_id = 6071 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 6072 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 6073 then
	sram_write <= x"820034A0";
end if;
if first_state_sram_input_id = 6074 then
	sram_write <= x"07DC0018";
end if;
if first_state_sram_input_id = 6075 then
	sram_write <= x"82005F10";
end if;
if first_state_sram_input_id = 6076 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 6077 then
	sram_write <= x"00460000";
end if;
if first_state_sram_input_id = 6078 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 6079 then
	sram_write <= x"03DC0018";
end if;
if first_state_sram_input_id = 6080 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 6081 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 6082 then
	sram_write <= x"820032A4";
end if;
if first_state_sram_input_id = 6083 then
	sram_write <= x"07DC0018";
end if;
if first_state_sram_input_id = 6084 then
	sram_write <= x"82005FF4";
end if;
if first_state_sram_input_id = 6085 then
	sram_write <= x"02C00000";
end if;
if first_state_sram_input_id = 6086 then
	sram_write <= x"02E00001";
end if;
if first_state_sram_input_id = 6087 then
	sram_write <= x"03000002";
end if;
if first_state_sram_input_id = 6088 then
	sram_write <= x"CC3C0010";
end if;
if first_state_sram_input_id = 6089 then
	sram_write <= x"CC7C0018";
end if;
if first_state_sram_input_id = 6090 then
	sram_write <= x"CC5C0020";
end if;
if first_state_sram_input_id = 6091 then
	sram_write <= x"C4BC0028";
end if;
if first_state_sram_input_id = 6092 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 6093 then
	sram_write <= x"008E0000";
end if;
if first_state_sram_input_id = 6094 then
	sram_write <= x"00460000";
end if;
if first_state_sram_input_id = 6095 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 6096 then
	sram_write <= x"00B00000";
end if;
if first_state_sram_input_id = 6097 then
	sram_write <= x"006C0000";
end if;
if first_state_sram_input_id = 6098 then
	sram_write <= x"03DC0034";
end if;
if first_state_sram_input_id = 6099 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 6100 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 6101 then
	sram_write <= x"8200317C";
end if;
if first_state_sram_input_id = 6102 then
	sram_write <= x"07DC0034";
end if;
if first_state_sram_input_id = 6103 then
	sram_write <= x"82205F68";
end if;
if first_state_sram_input_id = 6104 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 6105 then
	sram_write <= x"82005FF4";
end if;
if first_state_sram_input_id = 6106 then
	sram_write <= x"02600001";
end if;
if first_state_sram_input_id = 6107 then
	sram_write <= x"02800002";
end if;
if first_state_sram_input_id = 6108 then
	sram_write <= x"02A00000";
end if;
if first_state_sram_input_id = 6109 then
	sram_write <= x"C83C0020";
end if;
if first_state_sram_input_id = 6110 then
	sram_write <= x"C85C0018";
end if;
if first_state_sram_input_id = 6111 then
	sram_write <= x"C87C0010";
end if;
if first_state_sram_input_id = 6112 then
	sram_write <= x"C03C0028";
end if;
if first_state_sram_input_id = 6113 then
	sram_write <= x"C05C0000";
end if;
if first_state_sram_input_id = 6114 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 6115 then
	sram_write <= x"03DC0034";
end if;
if first_state_sram_input_id = 6116 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 6117 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 6118 then
	sram_write <= x"8200317C";
end if;
if first_state_sram_input_id = 6119 then
	sram_write <= x"07DC0034";
end if;
if first_state_sram_input_id = 6120 then
	sram_write <= x"82205FAC";
end if;
if first_state_sram_input_id = 6121 then
	sram_write <= x"02200002";
end if;
if first_state_sram_input_id = 6122 then
	sram_write <= x"82005FF4";
end if;
if first_state_sram_input_id = 6123 then
	sram_write <= x"02600002";
end if;
if first_state_sram_input_id = 6124 then
	sram_write <= x"02800000";
end if;
if first_state_sram_input_id = 6125 then
	sram_write <= x"02A00001";
end if;
if first_state_sram_input_id = 6126 then
	sram_write <= x"C83C0018";
end if;
if first_state_sram_input_id = 6127 then
	sram_write <= x"C85C0010";
end if;
if first_state_sram_input_id = 6128 then
	sram_write <= x"C87C0020";
end if;
if first_state_sram_input_id = 6129 then
	sram_write <= x"C03C0028";
end if;
if first_state_sram_input_id = 6130 then
	sram_write <= x"C05C0000";
end if;
if first_state_sram_input_id = 6131 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 6132 then
	sram_write <= x"03DC0034";
end if;
if first_state_sram_input_id = 6133 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 6134 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 6135 then
	sram_write <= x"8200317C";
end if;
if first_state_sram_input_id = 6136 then
	sram_write <= x"07DC0034";
end if;
if first_state_sram_input_id = 6137 then
	sram_write <= x"82205FF0";
end if;
if first_state_sram_input_id = 6138 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 6139 then
	sram_write <= x"82005FF4";
end if;
if first_state_sram_input_id = 6140 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 6141 then
	sram_write <= x"82206114";
end if;
if first_state_sram_input_id = 6142 then
	sram_write <= x"022002AC";
end if;
if first_state_sram_input_id = 6143 then
	sram_write <= x"C8220000";
end if;
if first_state_sram_input_id = 6144 then
	sram_write <= x"022002B4";
end if;
if first_state_sram_input_id = 6145 then
	sram_write <= x"C8420000";
end if;
if first_state_sram_input_id = 6146 then
	sram_write <= x"8E246010";
end if;
if first_state_sram_input_id = 6147 then
	sram_write <= x"82006110";
end if;
if first_state_sram_input_id = 6148 then
	sram_write <= x"C03C000C";
end if;
if first_state_sram_input_id = 6149 then
	sram_write <= x"C0420004";
end if;
if first_state_sram_input_id = 6150 then
	sram_write <= x"0260FFFF";
end if;
if first_state_sram_input_id = 6151 then
	sram_write <= x"82466110";
end if;
if first_state_sram_input_id = 6152 then
	sram_write <= x"026001E0";
end if;
if first_state_sram_input_id = 6153 then
	sram_write <= x"22440220";
end if;
if first_state_sram_input_id = 6154 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 6155 then
	sram_write <= x"02800000";
end if;
if first_state_sram_input_id = 6156 then
	sram_write <= x"C0BC0000";
end if;
if first_state_sram_input_id = 6157 then
	sram_write <= x"C47C002C";
end if;
if first_state_sram_input_id = 6158 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 6159 then
	sram_write <= x"006A0000";
end if;
if first_state_sram_input_id = 6160 then
	sram_write <= x"00280000";
end if;
if first_state_sram_input_id = 6161 then
	sram_write <= x"03DC0038";
end if;
if first_state_sram_input_id = 6162 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 6163 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 6164 then
	sram_write <= x"820057C8";
end if;
if first_state_sram_input_id = 6165 then
	sram_write <= x"07DC0038";
end if;
if first_state_sram_input_id = 6166 then
	sram_write <= x"C03C000C";
end if;
if first_state_sram_input_id = 6167 then
	sram_write <= x"C0420008";
end if;
if first_state_sram_input_id = 6168 then
	sram_write <= x"0260FFFF";
end if;
if first_state_sram_input_id = 6169 then
	sram_write <= x"8246610C";
end if;
if first_state_sram_input_id = 6170 then
	sram_write <= x"22440220";
end if;
if first_state_sram_input_id = 6171 then
	sram_write <= x"C07C002C";
end if;
if first_state_sram_input_id = 6172 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 6173 then
	sram_write <= x"02800000";
end if;
if first_state_sram_input_id = 6174 then
	sram_write <= x"C0BC0000";
end if;
if first_state_sram_input_id = 6175 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 6176 then
	sram_write <= x"006A0000";
end if;
if first_state_sram_input_id = 6177 then
	sram_write <= x"00280000";
end if;
if first_state_sram_input_id = 6178 then
	sram_write <= x"03DC0038";
end if;
if first_state_sram_input_id = 6179 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 6180 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 6181 then
	sram_write <= x"820057C8";
end if;
if first_state_sram_input_id = 6182 then
	sram_write <= x"07DC0038";
end if;
if first_state_sram_input_id = 6183 then
	sram_write <= x"C03C000C";
end if;
if first_state_sram_input_id = 6184 then
	sram_write <= x"C042000C";
end if;
if first_state_sram_input_id = 6185 then
	sram_write <= x"0260FFFF";
end if;
if first_state_sram_input_id = 6186 then
	sram_write <= x"82466108";
end if;
if first_state_sram_input_id = 6187 then
	sram_write <= x"22440220";
end if;
if first_state_sram_input_id = 6188 then
	sram_write <= x"C07C002C";
end if;
if first_state_sram_input_id = 6189 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 6190 then
	sram_write <= x"02600000";
end if;
if first_state_sram_input_id = 6191 then
	sram_write <= x"C09C0000";
end if;
if first_state_sram_input_id = 6192 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 6193 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 6194 then
	sram_write <= x"00680000";
end if;
if first_state_sram_input_id = 6195 then
	sram_write <= x"03DC0038";
end if;
if first_state_sram_input_id = 6196 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 6197 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 6198 then
	sram_write <= x"820057C8";
end if;
if first_state_sram_input_id = 6199 then
	sram_write <= x"07DC0038";
end if;
if first_state_sram_input_id = 6200 then
	sram_write <= x"02200004";
end if;
if first_state_sram_input_id = 6201 then
	sram_write <= x"C05C000C";
end if;
if first_state_sram_input_id = 6202 then
	sram_write <= x"C07C0000";
end if;
if first_state_sram_input_id = 6203 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 6204 then
	sram_write <= x"03DC0038";
end if;
if first_state_sram_input_id = 6205 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 6206 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 6207 then
	sram_write <= x"82005CDC";
end if;
if first_state_sram_input_id = 6208 then
	sram_write <= x"07DC0038";
end if;
if first_state_sram_input_id = 6209 then
	sram_write <= x"82006108";
end if;
if first_state_sram_input_id = 6210 then
	sram_write <= x"8200610C";
end if;
if first_state_sram_input_id = 6211 then
	sram_write <= x"82006110";
end if;
if first_state_sram_input_id = 6212 then
	sram_write <= x"82006114";
end if;
if first_state_sram_input_id = 6213 then
	sram_write <= x"82006214";
end if;
if first_state_sram_input_id = 6214 then
	sram_write <= x"C0A80004";
end if;
if first_state_sram_input_id = 6215 then
	sram_write <= x"02C0FFFF";
end if;
if first_state_sram_input_id = 6216 then
	sram_write <= x"82AC6214";
end if;
if first_state_sram_input_id = 6217 then
	sram_write <= x"02C001E0";
end if;
if first_state_sram_input_id = 6218 then
	sram_write <= x"22AA0220";
end if;
if first_state_sram_input_id = 6219 then
	sram_write <= x"D0ACA000";
end if;
if first_state_sram_input_id = 6220 then
	sram_write <= x"02E00000";
end if;
if first_state_sram_input_id = 6221 then
	sram_write <= x"C4DC0030";
end if;
if first_state_sram_input_id = 6222 then
	sram_write <= x"C49C000C";
end if;
if first_state_sram_input_id = 6223 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 6224 then
	sram_write <= x"004A0000";
end if;
if first_state_sram_input_id = 6225 then
	sram_write <= x"002E0000";
end if;
if first_state_sram_input_id = 6226 then
	sram_write <= x"03DC003C";
end if;
if first_state_sram_input_id = 6227 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 6228 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 6229 then
	sram_write <= x"820057C8";
end if;
if first_state_sram_input_id = 6230 then
	sram_write <= x"07DC003C";
end if;
if first_state_sram_input_id = 6231 then
	sram_write <= x"C03C000C";
end if;
if first_state_sram_input_id = 6232 then
	sram_write <= x"C0420008";
end if;
if first_state_sram_input_id = 6233 then
	sram_write <= x"0260FFFF";
end if;
if first_state_sram_input_id = 6234 then
	sram_write <= x"82466210";
end if;
if first_state_sram_input_id = 6235 then
	sram_write <= x"22440220";
end if;
if first_state_sram_input_id = 6236 then
	sram_write <= x"C07C0030";
end if;
if first_state_sram_input_id = 6237 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 6238 then
	sram_write <= x"02800000";
end if;
if first_state_sram_input_id = 6239 then
	sram_write <= x"C0BC0000";
end if;
if first_state_sram_input_id = 6240 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 6241 then
	sram_write <= x"006A0000";
end if;
if first_state_sram_input_id = 6242 then
	sram_write <= x"00280000";
end if;
if first_state_sram_input_id = 6243 then
	sram_write <= x"03DC003C";
end if;
if first_state_sram_input_id = 6244 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 6245 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 6246 then
	sram_write <= x"820057C8";
end if;
if first_state_sram_input_id = 6247 then
	sram_write <= x"07DC003C";
end if;
if first_state_sram_input_id = 6248 then
	sram_write <= x"C03C000C";
end if;
if first_state_sram_input_id = 6249 then
	sram_write <= x"C042000C";
end if;
if first_state_sram_input_id = 6250 then
	sram_write <= x"0260FFFF";
end if;
if first_state_sram_input_id = 6251 then
	sram_write <= x"8246620C";
end if;
if first_state_sram_input_id = 6252 then
	sram_write <= x"22440220";
end if;
if first_state_sram_input_id = 6253 then
	sram_write <= x"C07C0030";
end if;
if first_state_sram_input_id = 6254 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 6255 then
	sram_write <= x"02600000";
end if;
if first_state_sram_input_id = 6256 then
	sram_write <= x"C09C0000";
end if;
if first_state_sram_input_id = 6257 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 6258 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 6259 then
	sram_write <= x"00680000";
end if;
if first_state_sram_input_id = 6260 then
	sram_write <= x"03DC003C";
end if;
if first_state_sram_input_id = 6261 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 6262 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 6263 then
	sram_write <= x"820057C8";
end if;
if first_state_sram_input_id = 6264 then
	sram_write <= x"07DC003C";
end if;
if first_state_sram_input_id = 6265 then
	sram_write <= x"02200004";
end if;
if first_state_sram_input_id = 6266 then
	sram_write <= x"C05C000C";
end if;
if first_state_sram_input_id = 6267 then
	sram_write <= x"C07C0000";
end if;
if first_state_sram_input_id = 6268 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 6269 then
	sram_write <= x"03DC003C";
end if;
if first_state_sram_input_id = 6270 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 6271 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 6272 then
	sram_write <= x"82005CDC";
end if;
if first_state_sram_input_id = 6273 then
	sram_write <= x"07DC003C";
end if;
if first_state_sram_input_id = 6274 then
	sram_write <= x"8200620C";
end if;
if first_state_sram_input_id = 6275 then
	sram_write <= x"82006210";
end if;
if first_state_sram_input_id = 6276 then
	sram_write <= x"82006214";
end if;
if first_state_sram_input_id = 6277 then
	sram_write <= x"C03C0008";
end if;
if first_state_sram_input_id = 6278 then
	sram_write <= x"02220001";
end if;
if first_state_sram_input_id = 6279 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 6280 then
	sram_write <= x"C07C0004";
end if;
if first_state_sram_input_id = 6281 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 6282 then
	sram_write <= x"C0840000";
end if;
if first_state_sram_input_id = 6283 then
	sram_write <= x"02A0FFFF";
end if;
if first_state_sram_input_id = 6284 then
	sram_write <= x"828A641C";
end if;
if first_state_sram_input_id = 6285 then
	sram_write <= x"02A00063";
end if;
if first_state_sram_input_id = 6286 then
	sram_write <= x"C43C0034";
end if;
if first_state_sram_input_id = 6287 then
	sram_write <= x"828A634C";
end if;
if first_state_sram_input_id = 6288 then
	sram_write <= x"02A0030C";
end if;
if first_state_sram_input_id = 6289 then
	sram_write <= x"C0DC0000";
end if;
if first_state_sram_input_id = 6290 then
	sram_write <= x"C45C0038";
end if;
if first_state_sram_input_id = 6291 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 6292 then
	sram_write <= x"006A0000";
end if;
if first_state_sram_input_id = 6293 then
	sram_write <= x"004C0000";
end if;
if first_state_sram_input_id = 6294 then
	sram_write <= x"00280000";
end if;
if first_state_sram_input_id = 6295 then
	sram_write <= x"03DC0044";
end if;
if first_state_sram_input_id = 6296 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 6297 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 6298 then
	sram_write <= x"820036D4";
end if;
if first_state_sram_input_id = 6299 then
	sram_write <= x"07DC0044";
end if;
if first_state_sram_input_id = 6300 then
	sram_write <= x"82206348";
end if;
if first_state_sram_input_id = 6301 then
	sram_write <= x"022002AC";
end if;
if first_state_sram_input_id = 6302 then
	sram_write <= x"C8220000";
end if;
if first_state_sram_input_id = 6303 then
	sram_write <= x"022002B4";
end if;
if first_state_sram_input_id = 6304 then
	sram_write <= x"C8420000";
end if;
if first_state_sram_input_id = 6305 then
	sram_write <= x"8E24628C";
end if;
if first_state_sram_input_id = 6306 then
	sram_write <= x"82006344";
end if;
if first_state_sram_input_id = 6307 then
	sram_write <= x"C03C0038";
end if;
if first_state_sram_input_id = 6308 then
	sram_write <= x"C0420004";
end if;
if first_state_sram_input_id = 6309 then
	sram_write <= x"0260FFFF";
end if;
if first_state_sram_input_id = 6310 then
	sram_write <= x"82466344";
end if;
if first_state_sram_input_id = 6311 then
	sram_write <= x"026001E0";
end if;
if first_state_sram_input_id = 6312 then
	sram_write <= x"22440220";
end if;
if first_state_sram_input_id = 6313 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 6314 then
	sram_write <= x"02800000";
end if;
if first_state_sram_input_id = 6315 then
	sram_write <= x"C0BC0000";
end if;
if first_state_sram_input_id = 6316 then
	sram_write <= x"C47C003C";
end if;
if first_state_sram_input_id = 6317 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 6318 then
	sram_write <= x"006A0000";
end if;
if first_state_sram_input_id = 6319 then
	sram_write <= x"00280000";
end if;
if first_state_sram_input_id = 6320 then
	sram_write <= x"03DC0048";
end if;
if first_state_sram_input_id = 6321 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 6322 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 6323 then
	sram_write <= x"820057C8";
end if;
if first_state_sram_input_id = 6324 then
	sram_write <= x"07DC0048";
end if;
if first_state_sram_input_id = 6325 then
	sram_write <= x"C03C0038";
end if;
if first_state_sram_input_id = 6326 then
	sram_write <= x"C0420008";
end if;
if first_state_sram_input_id = 6327 then
	sram_write <= x"0260FFFF";
end if;
if first_state_sram_input_id = 6328 then
	sram_write <= x"82466340";
end if;
if first_state_sram_input_id = 6329 then
	sram_write <= x"22440220";
end if;
if first_state_sram_input_id = 6330 then
	sram_write <= x"C07C003C";
end if;
if first_state_sram_input_id = 6331 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 6332 then
	sram_write <= x"02600000";
end if;
if first_state_sram_input_id = 6333 then
	sram_write <= x"C09C0000";
end if;
if first_state_sram_input_id = 6334 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 6335 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 6336 then
	sram_write <= x"00680000";
end if;
if first_state_sram_input_id = 6337 then
	sram_write <= x"03DC0048";
end if;
if first_state_sram_input_id = 6338 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 6339 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 6340 then
	sram_write <= x"820057C8";
end if;
if first_state_sram_input_id = 6341 then
	sram_write <= x"07DC0048";
end if;
if first_state_sram_input_id = 6342 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 6343 then
	sram_write <= x"C05C0038";
end if;
if first_state_sram_input_id = 6344 then
	sram_write <= x"C07C0000";
end if;
if first_state_sram_input_id = 6345 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 6346 then
	sram_write <= x"03DC0048";
end if;
if first_state_sram_input_id = 6347 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 6348 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 6349 then
	sram_write <= x"82005CDC";
end if;
if first_state_sram_input_id = 6350 then
	sram_write <= x"07DC0048";
end if;
if first_state_sram_input_id = 6351 then
	sram_write <= x"82006340";
end if;
if first_state_sram_input_id = 6352 then
	sram_write <= x"82006344";
end if;
if first_state_sram_input_id = 6353 then
	sram_write <= x"82006348";
end if;
if first_state_sram_input_id = 6354 then
	sram_write <= x"82006408";
end if;
if first_state_sram_input_id = 6355 then
	sram_write <= x"C0840004";
end if;
if first_state_sram_input_id = 6356 then
	sram_write <= x"02A0FFFF";
end if;
if first_state_sram_input_id = 6357 then
	sram_write <= x"828A6408";
end if;
if first_state_sram_input_id = 6358 then
	sram_write <= x"02A001E0";
end if;
if first_state_sram_input_id = 6359 then
	sram_write <= x"22880220";
end if;
if first_state_sram_input_id = 6360 then
	sram_write <= x"D08A8000";
end if;
if first_state_sram_input_id = 6361 then
	sram_write <= x"02C00000";
end if;
if first_state_sram_input_id = 6362 then
	sram_write <= x"C0FC0000";
end if;
if first_state_sram_input_id = 6363 then
	sram_write <= x"C4BC0040";
end if;
if first_state_sram_input_id = 6364 then
	sram_write <= x"C45C0038";
end if;
if first_state_sram_input_id = 6365 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 6366 then
	sram_write <= x"006E0000";
end if;
if first_state_sram_input_id = 6367 then
	sram_write <= x"00480000";
end if;
if first_state_sram_input_id = 6368 then
	sram_write <= x"002C0000";
end if;
if first_state_sram_input_id = 6369 then
	sram_write <= x"03DC004C";
end if;
if first_state_sram_input_id = 6370 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 6371 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 6372 then
	sram_write <= x"820057C8";
end if;
if first_state_sram_input_id = 6373 then
	sram_write <= x"07DC004C";
end if;
if first_state_sram_input_id = 6374 then
	sram_write <= x"C03C0038";
end if;
if first_state_sram_input_id = 6375 then
	sram_write <= x"C0420008";
end if;
if first_state_sram_input_id = 6376 then
	sram_write <= x"0260FFFF";
end if;
if first_state_sram_input_id = 6377 then
	sram_write <= x"82466404";
end if;
if first_state_sram_input_id = 6378 then
	sram_write <= x"22440220";
end if;
if first_state_sram_input_id = 6379 then
	sram_write <= x"C07C0040";
end if;
if first_state_sram_input_id = 6380 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 6381 then
	sram_write <= x"02600000";
end if;
if first_state_sram_input_id = 6382 then
	sram_write <= x"C09C0000";
end if;
if first_state_sram_input_id = 6383 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 6384 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 6385 then
	sram_write <= x"00680000";
end if;
if first_state_sram_input_id = 6386 then
	sram_write <= x"03DC004C";
end if;
if first_state_sram_input_id = 6387 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 6388 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 6389 then
	sram_write <= x"820057C8";
end if;
if first_state_sram_input_id = 6390 then
	sram_write <= x"07DC004C";
end if;
if first_state_sram_input_id = 6391 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 6392 then
	sram_write <= x"C05C0038";
end if;
if first_state_sram_input_id = 6393 then
	sram_write <= x"C07C0000";
end if;
if first_state_sram_input_id = 6394 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 6395 then
	sram_write <= x"03DC004C";
end if;
if first_state_sram_input_id = 6396 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 6397 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 6398 then
	sram_write <= x"82005CDC";
end if;
if first_state_sram_input_id = 6399 then
	sram_write <= x"07DC004C";
end if;
if first_state_sram_input_id = 6400 then
	sram_write <= x"82006404";
end if;
if first_state_sram_input_id = 6401 then
	sram_write <= x"82006408";
end if;
if first_state_sram_input_id = 6402 then
	sram_write <= x"C03C0034";
end if;
if first_state_sram_input_id = 6403 then
	sram_write <= x"02220001";
end if;
if first_state_sram_input_id = 6404 then
	sram_write <= x"C05C0004";
end if;
if first_state_sram_input_id = 6405 then
	sram_write <= x"C07C0000";
end if;
if first_state_sram_input_id = 6406 then
	sram_write <= x"82005E4C";
end if;
if first_state_sram_input_id = 6407 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 6408 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 6409 then
	sram_write <= x"C0860000";
end if;
if first_state_sram_input_id = 6410 then
	sram_write <= x"22A20220";
end if;
if first_state_sram_input_id = 6411 then
	sram_write <= x"D0A4A000";
end if;
if first_state_sram_input_id = 6412 then
	sram_write <= x"02C0FFFF";
end if;
if first_state_sram_input_id = 6413 then
	sram_write <= x"82AC6874";
end if;
if first_state_sram_input_id = 6414 then
	sram_write <= x"02C000C8";
end if;
if first_state_sram_input_id = 6415 then
	sram_write <= x"22EA0220";
end if;
if first_state_sram_input_id = 6416 then
	sram_write <= x"D0ECE000";
end if;
if first_state_sram_input_id = 6417 then
	sram_write <= x"C10E0028";
end if;
if first_state_sram_input_id = 6418 then
	sram_write <= x"C8300000";
end if;
if first_state_sram_input_id = 6419 then
	sram_write <= x"C8500004";
end if;
if first_state_sram_input_id = 6420 then
	sram_write <= x"C8700008";
end if;
if first_state_sram_input_id = 6421 then
	sram_write <= x"C1260004";
end if;
if first_state_sram_input_id = 6422 then
	sram_write <= x"234A0220";
end if;
if first_state_sram_input_id = 6423 then
	sram_write <= x"D1334000";
end if;
if first_state_sram_input_id = 6424 then
	sram_write <= x"C14E0004";
end if;
if first_state_sram_input_id = 6425 then
	sram_write <= x"C49C0000";
end if;
if first_state_sram_input_id = 6426 then
	sram_write <= x"02800001";
end if;
if first_state_sram_input_id = 6427 then
	sram_write <= x"C47C0004";
end if;
if first_state_sram_input_id = 6428 then
	sram_write <= x"C45C0008";
end if;
if first_state_sram_input_id = 6429 then
	sram_write <= x"C43C000C";
end if;
if first_state_sram_input_id = 6430 then
	sram_write <= x"C4DC0010";
end if;
if first_state_sram_input_id = 6431 then
	sram_write <= x"C4BC0014";
end if;
if first_state_sram_input_id = 6432 then
	sram_write <= x"834864E0";
end if;
if first_state_sram_input_id = 6433 then
	sram_write <= x"02800002";
end if;
if first_state_sram_input_id = 6434 then
	sram_write <= x"834864B4";
end if;
if first_state_sram_input_id = 6435 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 6436 then
	sram_write <= x"00700000";
end if;
if first_state_sram_input_id = 6437 then
	sram_write <= x"00520000";
end if;
if first_state_sram_input_id = 6438 then
	sram_write <= x"002E0000";
end if;
if first_state_sram_input_id = 6439 then
	sram_write <= x"03DC0020";
end if;
if first_state_sram_input_id = 6440 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 6441 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 6442 then
	sram_write <= x"82003BD4";
end if;
if first_state_sram_input_id = 6443 then
	sram_write <= x"07DC0020";
end if;
if first_state_sram_input_id = 6444 then
	sram_write <= x"820064DC";
end if;
if first_state_sram_input_id = 6445 then
	sram_write <= x"C8320000";
end if;
if first_state_sram_input_id = 6446 then
	sram_write <= x"8E2064C4";
end if;
if first_state_sram_input_id = 6447 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 6448 then
	sram_write <= x"820064DC";
end if;
if first_state_sram_input_id = 6449 then
	sram_write <= x"028002AC";
end if;
if first_state_sram_input_id = 6450 then
	sram_write <= x"C8320000";
end if;
if first_state_sram_input_id = 6451 then
	sram_write <= x"C850000C";
end if;
if first_state_sram_input_id = 6452 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 6453 then
	sram_write <= x"CC280000";
end if;
if first_state_sram_input_id = 6454 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 6455 then
	sram_write <= x"82006508";
end if;
if first_state_sram_input_id = 6456 then
	sram_write <= x"C0860000";
end if;
if first_state_sram_input_id = 6457 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 6458 then
	sram_write <= x"00720000";
end if;
if first_state_sram_input_id = 6459 then
	sram_write <= x"00480000";
end if;
if first_state_sram_input_id = 6460 then
	sram_write <= x"002E0000";
end if;
if first_state_sram_input_id = 6461 then
	sram_write <= x"03DC0020";
end if;
if first_state_sram_input_id = 6462 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 6463 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 6464 then
	sram_write <= x"8200389C";
end if;
if first_state_sram_input_id = 6465 then
	sram_write <= x"07DC0020";
end if;
if first_state_sram_input_id = 6466 then
	sram_write <= x"82206844";
end if;
if first_state_sram_input_id = 6467 then
	sram_write <= x"024002AC";
end if;
if first_state_sram_input_id = 6468 then
	sram_write <= x"C8240000";
end if;
if first_state_sram_input_id = 6469 then
	sram_write <= x"8E02651C";
end if;
if first_state_sram_input_id = 6470 then
	sram_write <= x"82006830";
end if;
if first_state_sram_input_id = 6471 then
	sram_write <= x"024002B4";
end if;
if first_state_sram_input_id = 6472 then
	sram_write <= x"C8440000";
end if;
if first_state_sram_input_id = 6473 then
	sram_write <= x"8E24652C";
end if;
if first_state_sram_input_id = 6474 then
	sram_write <= x"82006830";
end if;
if first_state_sram_input_id = 6475 then
	sram_write <= x"C8400074";
end if;
if first_state_sram_input_id = 6476 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 6477 then
	sram_write <= x"C07C0000";
end if;
if first_state_sram_input_id = 6478 then
	sram_write <= x"C8460000";
end if;
if first_state_sram_input_id = 6479 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 6480 then
	sram_write <= x"02800318";
end if;
if first_state_sram_input_id = 6481 then
	sram_write <= x"C8680000";
end if;
if first_state_sram_input_id = 6482 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 6483 then
	sram_write <= x"C8660004";
end if;
if first_state_sram_input_id = 6484 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 6485 then
	sram_write <= x"C8880004";
end if;
if first_state_sram_input_id = 6486 then
	sram_write <= x"40668000";
end if;
if first_state_sram_input_id = 6487 then
	sram_write <= x"C8860008";
end if;
if first_state_sram_input_id = 6488 then
	sram_write <= x"48882000";
end if;
if first_state_sram_input_id = 6489 then
	sram_write <= x"C8A80008";
end if;
if first_state_sram_input_id = 6490 then
	sram_write <= x"4088A000";
end if;
if first_state_sram_input_id = 6491 then
	sram_write <= x"C07C0008";
end if;
if first_state_sram_input_id = 6492 then
	sram_write <= x"C0860000";
end if;
if first_state_sram_input_id = 6493 then
	sram_write <= x"02A0FFFF";
end if;
if first_state_sram_input_id = 6494 then
	sram_write <= x"C43C0018";
end if;
if first_state_sram_input_id = 6495 then
	sram_write <= x"CC9C0020";
end if;
if first_state_sram_input_id = 6496 then
	sram_write <= x"CC7C0028";
end if;
if first_state_sram_input_id = 6497 then
	sram_write <= x"CC5C0030";
end if;
if first_state_sram_input_id = 6498 then
	sram_write <= x"C45C0038";
end if;
if first_state_sram_input_id = 6499 then
	sram_write <= x"CC3C0040";
end if;
if first_state_sram_input_id = 6500 then
	sram_write <= x"828A67E4";
end if;
if first_state_sram_input_id = 6501 then
	sram_write <= x"22880220";
end if;
if first_state_sram_input_id = 6502 then
	sram_write <= x"C0BC0010";
end if;
if first_state_sram_input_id = 6503 then
	sram_write <= x"D08A8000";
end if;
if first_state_sram_input_id = 6504 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 6505 then
	sram_write <= x"00280000";
end if;
if first_state_sram_input_id = 6506 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 6507 then
	sram_write <= x"40406000";
end if;
if first_state_sram_input_id = 6508 then
	sram_write <= x"40608000";
end if;
if first_state_sram_input_id = 6509 then
	sram_write <= x"03DC0050";
end if;
if first_state_sram_input_id = 6510 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 6511 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 6512 then
	sram_write <= x"82004860";
end if;
if first_state_sram_input_id = 6513 then
	sram_write <= x"07DC0050";
end if;
if first_state_sram_input_id = 6514 then
	sram_write <= x"822065D4";
end if;
if first_state_sram_input_id = 6515 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 6516 then
	sram_write <= x"820067E0";
end if;
if first_state_sram_input_id = 6517 then
	sram_write <= x"C05C0008";
end if;
if first_state_sram_input_id = 6518 then
	sram_write <= x"C0240004";
end if;
if first_state_sram_input_id = 6519 then
	sram_write <= x"0260FFFF";
end if;
if first_state_sram_input_id = 6520 then
	sram_write <= x"822667DC";
end if;
if first_state_sram_input_id = 6521 then
	sram_write <= x"22220220";
end if;
if first_state_sram_input_id = 6522 then
	sram_write <= x"C07C0010";
end if;
if first_state_sram_input_id = 6523 then
	sram_write <= x"D0262000";
end if;
if first_state_sram_input_id = 6524 then
	sram_write <= x"C0820014";
end if;
if first_state_sram_input_id = 6525 then
	sram_write <= x"C8280000";
end if;
if first_state_sram_input_id = 6526 then
	sram_write <= x"C85C0030";
end if;
if first_state_sram_input_id = 6527 then
	sram_write <= x"44242000";
end if;
if first_state_sram_input_id = 6528 then
	sram_write <= x"C0820014";
end if;
if first_state_sram_input_id = 6529 then
	sram_write <= x"C8680004";
end if;
if first_state_sram_input_id = 6530 then
	sram_write <= x"C89C0028";
end if;
if first_state_sram_input_id = 6531 then
	sram_write <= x"44686000";
end if;
if first_state_sram_input_id = 6532 then
	sram_write <= x"C0820014";
end if;
if first_state_sram_input_id = 6533 then
	sram_write <= x"C8A80008";
end if;
if first_state_sram_input_id = 6534 then
	sram_write <= x"C8DC0020";
end if;
if first_state_sram_input_id = 6535 then
	sram_write <= x"44ACA000";
end if;
if first_state_sram_input_id = 6536 then
	sram_write <= x"C0820004";
end if;
if first_state_sram_input_id = 6537 then
	sram_write <= x"02A00001";
end if;
if first_state_sram_input_id = 6538 then
	sram_write <= x"828A66C0";
end if;
if first_state_sram_input_id = 6539 then
	sram_write <= x"02A00002";
end if;
if first_state_sram_input_id = 6540 then
	sram_write <= x"828A6658";
end if;
if first_state_sram_input_id = 6541 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 6542 then
	sram_write <= x"40406000";
end if;
if first_state_sram_input_id = 6543 then
	sram_write <= x"4060A000";
end if;
if first_state_sram_input_id = 6544 then
	sram_write <= x"03DC0050";
end if;
if first_state_sram_input_id = 6545 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 6546 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 6547 then
	sram_write <= x"82004780";
end if;
if first_state_sram_input_id = 6548 then
	sram_write <= x"07DC0050";
end if;
if first_state_sram_input_id = 6549 then
	sram_write <= x"820066BC";
end if;
if first_state_sram_input_id = 6550 then
	sram_write <= x"C0820010";
end if;
if first_state_sram_input_id = 6551 then
	sram_write <= x"C8E80000";
end if;
if first_state_sram_input_id = 6552 then
	sram_write <= x"482E2000";
end if;
if first_state_sram_input_id = 6553 then
	sram_write <= x"C8E80004";
end if;
if first_state_sram_input_id = 6554 then
	sram_write <= x"486E6000";
end if;
if first_state_sram_input_id = 6555 then
	sram_write <= x"40226000";
end if;
if first_state_sram_input_id = 6556 then
	sram_write <= x"C8680008";
end if;
if first_state_sram_input_id = 6557 then
	sram_write <= x"4866A000";
end if;
if first_state_sram_input_id = 6558 then
	sram_write <= x"40226000";
end if;
if first_state_sram_input_id = 6559 then
	sram_write <= x"C0220018";
end if;
if first_state_sram_input_id = 6560 then
	sram_write <= x"8E20668C";
end if;
if first_state_sram_input_id = 6561 then
	sram_write <= x"02800000";
end if;
if first_state_sram_input_id = 6562 then
	sram_write <= x"82006690";
end if;
if first_state_sram_input_id = 6563 then
	sram_write <= x"02800001";
end if;
if first_state_sram_input_id = 6564 then
	sram_write <= x"822066A8";
end if;
if first_state_sram_input_id = 6565 then
	sram_write <= x"8E2066A0";
end if;
if first_state_sram_input_id = 6566 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 6567 then
	sram_write <= x"820066A4";
end if;
if first_state_sram_input_id = 6568 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 6569 then
	sram_write <= x"820066AC";
end if;
if first_state_sram_input_id = 6570 then
	sram_write <= x"00280000";
end if;
if first_state_sram_input_id = 6571 then
	sram_write <= x"822066B8";
end if;
if first_state_sram_input_id = 6572 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 6573 then
	sram_write <= x"820066BC";
end if;
if first_state_sram_input_id = 6574 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 6575 then
	sram_write <= x"8200674C";
end if;
if first_state_sram_input_id = 6576 then
	sram_write <= x"8E2066C8";
end if;
if first_state_sram_input_id = 6577 then
	sram_write <= x"820066CC";
end if;
if first_state_sram_input_id = 6578 then
	sram_write <= x"44202000";
end if;
if first_state_sram_input_id = 6579 then
	sram_write <= x"C0820010";
end if;
if first_state_sram_input_id = 6580 then
	sram_write <= x"C8E80000";
end if;
if first_state_sram_input_id = 6581 then
	sram_write <= x"8E2E66E0";
end if;
if first_state_sram_input_id = 6582 then
	sram_write <= x"02800000";
end if;
if first_state_sram_input_id = 6583 then
	sram_write <= x"8200672C";
end if;
if first_state_sram_input_id = 6584 then
	sram_write <= x"8E6066EC";
end if;
if first_state_sram_input_id = 6585 then
	sram_write <= x"40206000";
end if;
if first_state_sram_input_id = 6586 then
	sram_write <= x"820066F0";
end if;
if first_state_sram_input_id = 6587 then
	sram_write <= x"44206000";
end if;
if first_state_sram_input_id = 6588 then
	sram_write <= x"C0820010";
end if;
if first_state_sram_input_id = 6589 then
	sram_write <= x"C8680004";
end if;
if first_state_sram_input_id = 6590 then
	sram_write <= x"8E266704";
end if;
if first_state_sram_input_id = 6591 then
	sram_write <= x"02800000";
end if;
if first_state_sram_input_id = 6592 then
	sram_write <= x"8200672C";
end if;
if first_state_sram_input_id = 6593 then
	sram_write <= x"8EA06710";
end if;
if first_state_sram_input_id = 6594 then
	sram_write <= x"4020A000";
end if;
if first_state_sram_input_id = 6595 then
	sram_write <= x"82006714";
end if;
if first_state_sram_input_id = 6596 then
	sram_write <= x"4420A000";
end if;
if first_state_sram_input_id = 6597 then
	sram_write <= x"C0820010";
end if;
if first_state_sram_input_id = 6598 then
	sram_write <= x"C8680008";
end if;
if first_state_sram_input_id = 6599 then
	sram_write <= x"8E266728";
end if;
if first_state_sram_input_id = 6600 then
	sram_write <= x"02800000";
end if;
if first_state_sram_input_id = 6601 then
	sram_write <= x"8200672C";
end if;
if first_state_sram_input_id = 6602 then
	sram_write <= x"02800001";
end if;
if first_state_sram_input_id = 6603 then
	sram_write <= x"82806738";
end if;
if first_state_sram_input_id = 6604 then
	sram_write <= x"C0220018";
end if;
if first_state_sram_input_id = 6605 then
	sram_write <= x"8200674C";
end if;
if first_state_sram_input_id = 6606 then
	sram_write <= x"C0220018";
end if;
if first_state_sram_input_id = 6607 then
	sram_write <= x"82206748";
end if;
if first_state_sram_input_id = 6608 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 6609 then
	sram_write <= x"8200674C";
end if;
if first_state_sram_input_id = 6610 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 6611 then
	sram_write <= x"82206758";
end if;
if first_state_sram_input_id = 6612 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 6613 then
	sram_write <= x"820067D8";
end if;
if first_state_sram_input_id = 6614 then
	sram_write <= x"C05C0008";
end if;
if first_state_sram_input_id = 6615 then
	sram_write <= x"C0240008";
end if;
if first_state_sram_input_id = 6616 then
	sram_write <= x"0260FFFF";
end if;
if first_state_sram_input_id = 6617 then
	sram_write <= x"822667D4";
end if;
if first_state_sram_input_id = 6618 then
	sram_write <= x"22220220";
end if;
if first_state_sram_input_id = 6619 then
	sram_write <= x"C07C0010";
end if;
if first_state_sram_input_id = 6620 then
	sram_write <= x"D0262000";
end if;
if first_state_sram_input_id = 6621 then
	sram_write <= x"C83C0030";
end if;
if first_state_sram_input_id = 6622 then
	sram_write <= x"C85C0028";
end if;
if first_state_sram_input_id = 6623 then
	sram_write <= x"C87C0020";
end if;
if first_state_sram_input_id = 6624 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 6625 then
	sram_write <= x"03DC0050";
end if;
if first_state_sram_input_id = 6626 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 6627 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 6628 then
	sram_write <= x"82004860";
end if;
if first_state_sram_input_id = 6629 then
	sram_write <= x"07DC0050";
end if;
if first_state_sram_input_id = 6630 then
	sram_write <= x"822067A4";
end if;
if first_state_sram_input_id = 6631 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 6632 then
	sram_write <= x"820067D0";
end if;
if first_state_sram_input_id = 6633 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 6634 then
	sram_write <= x"C83C0030";
end if;
if first_state_sram_input_id = 6635 then
	sram_write <= x"C85C0028";
end if;
if first_state_sram_input_id = 6636 then
	sram_write <= x"C87C0020";
end if;
if first_state_sram_input_id = 6637 then
	sram_write <= x"C05C0008";
end if;
if first_state_sram_input_id = 6638 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 6639 then
	sram_write <= x"03DC0050";
end if;
if first_state_sram_input_id = 6640 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 6641 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 6642 then
	sram_write <= x"82004A0C";
end if;
if first_state_sram_input_id = 6643 then
	sram_write <= x"07DC0050";
end if;
if first_state_sram_input_id = 6644 then
	sram_write <= x"820067D8";
end if;
if first_state_sram_input_id = 6645 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 6646 then
	sram_write <= x"820067E0";
end if;
if first_state_sram_input_id = 6647 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 6648 then
	sram_write <= x"820067E8";
end if;
if first_state_sram_input_id = 6649 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 6650 then
	sram_write <= x"82206830";
end if;
if first_state_sram_input_id = 6651 then
	sram_write <= x"C03C0038";
end if;
if first_state_sram_input_id = 6652 then
	sram_write <= x"C83C0040";
end if;
if first_state_sram_input_id = 6653 then
	sram_write <= x"CC220000";
end if;
if first_state_sram_input_id = 6654 then
	sram_write <= x"022002B8";
end if;
if first_state_sram_input_id = 6655 then
	sram_write <= x"C83C0030";
end if;
if first_state_sram_input_id = 6656 then
	sram_write <= x"CC220000";
end if;
if first_state_sram_input_id = 6657 then
	sram_write <= x"C83C0028";
end if;
if first_state_sram_input_id = 6658 then
	sram_write <= x"CC220004";
end if;
if first_state_sram_input_id = 6659 then
	sram_write <= x"C83C0020";
end if;
if first_state_sram_input_id = 6660 then
	sram_write <= x"CC220008";
end if;
if first_state_sram_input_id = 6661 then
	sram_write <= x"022002C4";
end if;
if first_state_sram_input_id = 6662 then
	sram_write <= x"C05C0014";
end if;
if first_state_sram_input_id = 6663 then
	sram_write <= x"C4420000";
end if;
if first_state_sram_input_id = 6664 then
	sram_write <= x"022002B0";
end if;
if first_state_sram_input_id = 6665 then
	sram_write <= x"C05C0018";
end if;
if first_state_sram_input_id = 6666 then
	sram_write <= x"C4420000";
end if;
if first_state_sram_input_id = 6667 then
	sram_write <= x"82006830";
end if;
if first_state_sram_input_id = 6668 then
	sram_write <= x"C03C000C";
end if;
if first_state_sram_input_id = 6669 then
	sram_write <= x"02220001";
end if;
if first_state_sram_input_id = 6670 then
	sram_write <= x"C05C0008";
end if;
if first_state_sram_input_id = 6671 then
	sram_write <= x"C07C0004";
end if;
if first_state_sram_input_id = 6672 then
	sram_write <= x"82006424";
end if;
if first_state_sram_input_id = 6673 then
	sram_write <= x"C03C0014";
end if;
if first_state_sram_input_id = 6674 then
	sram_write <= x"22220220";
end if;
if first_state_sram_input_id = 6675 then
	sram_write <= x"C05C0010";
end if;
if first_state_sram_input_id = 6676 then
	sram_write <= x"D0242000";
end if;
if first_state_sram_input_id = 6677 then
	sram_write <= x"C0220018";
end if;
if first_state_sram_input_id = 6678 then
	sram_write <= x"82206870";
end if;
if first_state_sram_input_id = 6679 then
	sram_write <= x"C03C000C";
end if;
if first_state_sram_input_id = 6680 then
	sram_write <= x"02220001";
end if;
if first_state_sram_input_id = 6681 then
	sram_write <= x"C05C0008";
end if;
if first_state_sram_input_id = 6682 then
	sram_write <= x"C07C0004";
end if;
if first_state_sram_input_id = 6683 then
	sram_write <= x"82006424";
end if;
if first_state_sram_input_id = 6684 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 6685 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 6686 then
	sram_write <= x"22820220";
end if;
if first_state_sram_input_id = 6687 then
	sram_write <= x"D0848000";
end if;
if first_state_sram_input_id = 6688 then
	sram_write <= x"02A0FFFF";
end if;
if first_state_sram_input_id = 6689 then
	sram_write <= x"828A69E4";
end if;
if first_state_sram_input_id = 6690 then
	sram_write <= x"02A001E0";
end if;
if first_state_sram_input_id = 6691 then
	sram_write <= x"22880220";
end if;
if first_state_sram_input_id = 6692 then
	sram_write <= x"D08A8000";
end if;
if first_state_sram_input_id = 6693 then
	sram_write <= x"02C00000";
end if;
if first_state_sram_input_id = 6694 then
	sram_write <= x"C47C0000";
end if;
if first_state_sram_input_id = 6695 then
	sram_write <= x"C4BC0004";
end if;
if first_state_sram_input_id = 6696 then
	sram_write <= x"C45C0008";
end if;
if first_state_sram_input_id = 6697 then
	sram_write <= x"C43C000C";
end if;
if first_state_sram_input_id = 6698 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 6699 then
	sram_write <= x"00480000";
end if;
if first_state_sram_input_id = 6700 then
	sram_write <= x"002C0000";
end if;
if first_state_sram_input_id = 6701 then
	sram_write <= x"03DC0018";
end if;
if first_state_sram_input_id = 6702 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 6703 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 6704 then
	sram_write <= x"82006424";
end if;
if first_state_sram_input_id = 6705 then
	sram_write <= x"07DC0018";
end if;
if first_state_sram_input_id = 6706 then
	sram_write <= x"C03C000C";
end if;
if first_state_sram_input_id = 6707 then
	sram_write <= x"02220001";
end if;
if first_state_sram_input_id = 6708 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 6709 then
	sram_write <= x"C07C0008";
end if;
if first_state_sram_input_id = 6710 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 6711 then
	sram_write <= x"0280FFFF";
end if;
if first_state_sram_input_id = 6712 then
	sram_write <= x"824869E0";
end if;
if first_state_sram_input_id = 6713 then
	sram_write <= x"22440220";
end if;
if first_state_sram_input_id = 6714 then
	sram_write <= x"C09C0004";
end if;
if first_state_sram_input_id = 6715 then
	sram_write <= x"D0484000";
end if;
if first_state_sram_input_id = 6716 then
	sram_write <= x"02A00000";
end if;
if first_state_sram_input_id = 6717 then
	sram_write <= x"C0DC0000";
end if;
if first_state_sram_input_id = 6718 then
	sram_write <= x"C43C0010";
end if;
if first_state_sram_input_id = 6719 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 6720 then
	sram_write <= x"006C0000";
end if;
if first_state_sram_input_id = 6721 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 6722 then
	sram_write <= x"03DC001C";
end if;
if first_state_sram_input_id = 6723 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 6724 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 6725 then
	sram_write <= x"82006424";
end if;
if first_state_sram_input_id = 6726 then
	sram_write <= x"07DC001C";
end if;
if first_state_sram_input_id = 6727 then
	sram_write <= x"C03C0010";
end if;
if first_state_sram_input_id = 6728 then
	sram_write <= x"02220001";
end if;
if first_state_sram_input_id = 6729 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 6730 then
	sram_write <= x"C07C0008";
end if;
if first_state_sram_input_id = 6731 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 6732 then
	sram_write <= x"0280FFFF";
end if;
if first_state_sram_input_id = 6733 then
	sram_write <= x"824869DC";
end if;
if first_state_sram_input_id = 6734 then
	sram_write <= x"22440220";
end if;
if first_state_sram_input_id = 6735 then
	sram_write <= x"C09C0004";
end if;
if first_state_sram_input_id = 6736 then
	sram_write <= x"D0484000";
end if;
if first_state_sram_input_id = 6737 then
	sram_write <= x"02A00000";
end if;
if first_state_sram_input_id = 6738 then
	sram_write <= x"C0DC0000";
end if;
if first_state_sram_input_id = 6739 then
	sram_write <= x"C43C0014";
end if;
if first_state_sram_input_id = 6740 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 6741 then
	sram_write <= x"006C0000";
end if;
if first_state_sram_input_id = 6742 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 6743 then
	sram_write <= x"03DC0020";
end if;
if first_state_sram_input_id = 6744 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 6745 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 6746 then
	sram_write <= x"82006424";
end if;
if first_state_sram_input_id = 6747 then
	sram_write <= x"07DC0020";
end if;
if first_state_sram_input_id = 6748 then
	sram_write <= x"C03C0014";
end if;
if first_state_sram_input_id = 6749 then
	sram_write <= x"02220001";
end if;
if first_state_sram_input_id = 6750 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 6751 then
	sram_write <= x"C07C0008";
end if;
if first_state_sram_input_id = 6752 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 6753 then
	sram_write <= x"0280FFFF";
end if;
if first_state_sram_input_id = 6754 then
	sram_write <= x"824869D8";
end if;
if first_state_sram_input_id = 6755 then
	sram_write <= x"22440220";
end if;
if first_state_sram_input_id = 6756 then
	sram_write <= x"C09C0004";
end if;
if first_state_sram_input_id = 6757 then
	sram_write <= x"D0484000";
end if;
if first_state_sram_input_id = 6758 then
	sram_write <= x"02800000";
end if;
if first_state_sram_input_id = 6759 then
	sram_write <= x"C0BC0000";
end if;
if first_state_sram_input_id = 6760 then
	sram_write <= x"C43C0018";
end if;
if first_state_sram_input_id = 6761 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 6762 then
	sram_write <= x"006A0000";
end if;
if first_state_sram_input_id = 6763 then
	sram_write <= x"00280000";
end if;
if first_state_sram_input_id = 6764 then
	sram_write <= x"03DC0024";
end if;
if first_state_sram_input_id = 6765 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 6766 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 6767 then
	sram_write <= x"82006424";
end if;
if first_state_sram_input_id = 6768 then
	sram_write <= x"07DC0024";
end if;
if first_state_sram_input_id = 6769 then
	sram_write <= x"C03C0018";
end if;
if first_state_sram_input_id = 6770 then
	sram_write <= x"02220001";
end if;
if first_state_sram_input_id = 6771 then
	sram_write <= x"C05C0008";
end if;
if first_state_sram_input_id = 6772 then
	sram_write <= x"C07C0000";
end if;
if first_state_sram_input_id = 6773 then
	sram_write <= x"82006878";
end if;
if first_state_sram_input_id = 6774 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 6775 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 6776 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 6777 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 6778 then
	sram_write <= x"22820220";
end if;
if first_state_sram_input_id = 6779 then
	sram_write <= x"D0848000";
end if;
if first_state_sram_input_id = 6780 then
	sram_write <= x"C0A80000";
end if;
if first_state_sram_input_id = 6781 then
	sram_write <= x"02C0FFFF";
end if;
if first_state_sram_input_id = 6782 then
	sram_write <= x"82AC6F88";
end if;
if first_state_sram_input_id = 6783 then
	sram_write <= x"02C00063";
end if;
if first_state_sram_input_id = 6784 then
	sram_write <= x"C47C0000";
end if;
if first_state_sram_input_id = 6785 then
	sram_write <= x"C45C0004";
end if;
if first_state_sram_input_id = 6786 then
	sram_write <= x"C43C0008";
end if;
if first_state_sram_input_id = 6787 then
	sram_write <= x"82AC6BF0";
end if;
if first_state_sram_input_id = 6788 then
	sram_write <= x"02C000C8";
end if;
if first_state_sram_input_id = 6789 then
	sram_write <= x"22EA0220";
end if;
if first_state_sram_input_id = 6790 then
	sram_write <= x"D0CCE000";
end if;
if first_state_sram_input_id = 6791 then
	sram_write <= x"C0EC0028";
end if;
if first_state_sram_input_id = 6792 then
	sram_write <= x"C82E0000";
end if;
if first_state_sram_input_id = 6793 then
	sram_write <= x"C84E0004";
end if;
if first_state_sram_input_id = 6794 then
	sram_write <= x"C86E0008";
end if;
if first_state_sram_input_id = 6795 then
	sram_write <= x"C1060004";
end if;
if first_state_sram_input_id = 6796 then
	sram_write <= x"22AA0220";
end if;
if first_state_sram_input_id = 6797 then
	sram_write <= x"D0B0A000";
end if;
if first_state_sram_input_id = 6798 then
	sram_write <= x"C10C0004";
end if;
if first_state_sram_input_id = 6799 then
	sram_write <= x"03200001";
end if;
if first_state_sram_input_id = 6800 then
	sram_write <= x"C49C000C";
end if;
if first_state_sram_input_id = 6801 then
	sram_write <= x"83126AA4";
end if;
if first_state_sram_input_id = 6802 then
	sram_write <= x"03200002";
end if;
if first_state_sram_input_id = 6803 then
	sram_write <= x"83126A78";
end if;
if first_state_sram_input_id = 6804 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 6805 then
	sram_write <= x"006E0000";
end if;
if first_state_sram_input_id = 6806 then
	sram_write <= x"004A0000";
end if;
if first_state_sram_input_id = 6807 then
	sram_write <= x"002C0000";
end if;
if first_state_sram_input_id = 6808 then
	sram_write <= x"03DC0018";
end if;
if first_state_sram_input_id = 6809 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 6810 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 6811 then
	sram_write <= x"82003BD4";
end if;
if first_state_sram_input_id = 6812 then
	sram_write <= x"07DC0018";
end if;
if first_state_sram_input_id = 6813 then
	sram_write <= x"82006AA0";
end if;
if first_state_sram_input_id = 6814 then
	sram_write <= x"C82A0000";
end if;
if first_state_sram_input_id = 6815 then
	sram_write <= x"8E206A88";
end if;
if first_state_sram_input_id = 6816 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 6817 then
	sram_write <= x"82006AA0";
end if;
if first_state_sram_input_id = 6818 then
	sram_write <= x"02C002AC";
end if;
if first_state_sram_input_id = 6819 then
	sram_write <= x"C82A0000";
end if;
if first_state_sram_input_id = 6820 then
	sram_write <= x"C84E000C";
end if;
if first_state_sram_input_id = 6821 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 6822 then
	sram_write <= x"CC2C0000";
end if;
if first_state_sram_input_id = 6823 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 6824 then
	sram_write <= x"82006ACC";
end if;
if first_state_sram_input_id = 6825 then
	sram_write <= x"C0E60000";
end if;
if first_state_sram_input_id = 6826 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 6827 then
	sram_write <= x"006A0000";
end if;
if first_state_sram_input_id = 6828 then
	sram_write <= x"004E0000";
end if;
if first_state_sram_input_id = 6829 then
	sram_write <= x"002C0000";
end if;
if first_state_sram_input_id = 6830 then
	sram_write <= x"03DC0018";
end if;
if first_state_sram_input_id = 6831 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 6832 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 6833 then
	sram_write <= x"8200389C";
end if;
if first_state_sram_input_id = 6834 then
	sram_write <= x"07DC0018";
end if;
if first_state_sram_input_id = 6835 then
	sram_write <= x"82206BEC";
end if;
if first_state_sram_input_id = 6836 then
	sram_write <= x"022002AC";
end if;
if first_state_sram_input_id = 6837 then
	sram_write <= x"C8220000";
end if;
if first_state_sram_input_id = 6838 then
	sram_write <= x"022002B4";
end if;
if first_state_sram_input_id = 6839 then
	sram_write <= x"C8420000";
end if;
if first_state_sram_input_id = 6840 then
	sram_write <= x"8E246AE8";
end if;
if first_state_sram_input_id = 6841 then
	sram_write <= x"82006BE8";
end if;
if first_state_sram_input_id = 6842 then
	sram_write <= x"C03C000C";
end if;
if first_state_sram_input_id = 6843 then
	sram_write <= x"C0420004";
end if;
if first_state_sram_input_id = 6844 then
	sram_write <= x"0260FFFF";
end if;
if first_state_sram_input_id = 6845 then
	sram_write <= x"82466BE8";
end if;
if first_state_sram_input_id = 6846 then
	sram_write <= x"026001E0";
end if;
if first_state_sram_input_id = 6847 then
	sram_write <= x"22440220";
end if;
if first_state_sram_input_id = 6848 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 6849 then
	sram_write <= x"02800000";
end if;
if first_state_sram_input_id = 6850 then
	sram_write <= x"C0BC0000";
end if;
if first_state_sram_input_id = 6851 then
	sram_write <= x"C47C0010";
end if;
if first_state_sram_input_id = 6852 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 6853 then
	sram_write <= x"006A0000";
end if;
if first_state_sram_input_id = 6854 then
	sram_write <= x"00280000";
end if;
if first_state_sram_input_id = 6855 then
	sram_write <= x"03DC001C";
end if;
if first_state_sram_input_id = 6856 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 6857 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 6858 then
	sram_write <= x"82006424";
end if;
if first_state_sram_input_id = 6859 then
	sram_write <= x"07DC001C";
end if;
if first_state_sram_input_id = 6860 then
	sram_write <= x"C03C000C";
end if;
if first_state_sram_input_id = 6861 then
	sram_write <= x"C0420008";
end if;
if first_state_sram_input_id = 6862 then
	sram_write <= x"0260FFFF";
end if;
if first_state_sram_input_id = 6863 then
	sram_write <= x"82466BE4";
end if;
if first_state_sram_input_id = 6864 then
	sram_write <= x"22440220";
end if;
if first_state_sram_input_id = 6865 then
	sram_write <= x"C07C0010";
end if;
if first_state_sram_input_id = 6866 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 6867 then
	sram_write <= x"02800000";
end if;
if first_state_sram_input_id = 6868 then
	sram_write <= x"C0BC0000";
end if;
if first_state_sram_input_id = 6869 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 6870 then
	sram_write <= x"006A0000";
end if;
if first_state_sram_input_id = 6871 then
	sram_write <= x"00280000";
end if;
if first_state_sram_input_id = 6872 then
	sram_write <= x"03DC001C";
end if;
if first_state_sram_input_id = 6873 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 6874 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 6875 then
	sram_write <= x"82006424";
end if;
if first_state_sram_input_id = 6876 then
	sram_write <= x"07DC001C";
end if;
if first_state_sram_input_id = 6877 then
	sram_write <= x"C03C000C";
end if;
if first_state_sram_input_id = 6878 then
	sram_write <= x"C042000C";
end if;
if first_state_sram_input_id = 6879 then
	sram_write <= x"0260FFFF";
end if;
if first_state_sram_input_id = 6880 then
	sram_write <= x"82466BE0";
end if;
if first_state_sram_input_id = 6881 then
	sram_write <= x"22440220";
end if;
if first_state_sram_input_id = 6882 then
	sram_write <= x"C07C0010";
end if;
if first_state_sram_input_id = 6883 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 6884 then
	sram_write <= x"02600000";
end if;
if first_state_sram_input_id = 6885 then
	sram_write <= x"C09C0000";
end if;
if first_state_sram_input_id = 6886 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 6887 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 6888 then
	sram_write <= x"00680000";
end if;
if first_state_sram_input_id = 6889 then
	sram_write <= x"03DC001C";
end if;
if first_state_sram_input_id = 6890 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 6891 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 6892 then
	sram_write <= x"82006424";
end if;
if first_state_sram_input_id = 6893 then
	sram_write <= x"07DC001C";
end if;
if first_state_sram_input_id = 6894 then
	sram_write <= x"02200004";
end if;
if first_state_sram_input_id = 6895 then
	sram_write <= x"C05C000C";
end if;
if first_state_sram_input_id = 6896 then
	sram_write <= x"C07C0000";
end if;
if first_state_sram_input_id = 6897 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 6898 then
	sram_write <= x"03DC001C";
end if;
if first_state_sram_input_id = 6899 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 6900 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 6901 then
	sram_write <= x"82006878";
end if;
if first_state_sram_input_id = 6902 then
	sram_write <= x"07DC001C";
end if;
if first_state_sram_input_id = 6903 then
	sram_write <= x"82006BE0";
end if;
if first_state_sram_input_id = 6904 then
	sram_write <= x"82006BE4";
end if;
if first_state_sram_input_id = 6905 then
	sram_write <= x"82006BE8";
end if;
if first_state_sram_input_id = 6906 then
	sram_write <= x"82006BEC";
end if;
if first_state_sram_input_id = 6907 then
	sram_write <= x"82006CEC";
end if;
if first_state_sram_input_id = 6908 then
	sram_write <= x"C0A80004";
end if;
if first_state_sram_input_id = 6909 then
	sram_write <= x"02C0FFFF";
end if;
if first_state_sram_input_id = 6910 then
	sram_write <= x"82AC6CEC";
end if;
if first_state_sram_input_id = 6911 then
	sram_write <= x"02C001E0";
end if;
if first_state_sram_input_id = 6912 then
	sram_write <= x"22AA0220";
end if;
if first_state_sram_input_id = 6913 then
	sram_write <= x"D0ACA000";
end if;
if first_state_sram_input_id = 6914 then
	sram_write <= x"02E00000";
end if;
if first_state_sram_input_id = 6915 then
	sram_write <= x"C4DC0014";
end if;
if first_state_sram_input_id = 6916 then
	sram_write <= x"C49C000C";
end if;
if first_state_sram_input_id = 6917 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 6918 then
	sram_write <= x"004A0000";
end if;
if first_state_sram_input_id = 6919 then
	sram_write <= x"002E0000";
end if;
if first_state_sram_input_id = 6920 then
	sram_write <= x"03DC0020";
end if;
if first_state_sram_input_id = 6921 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 6922 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 6923 then
	sram_write <= x"82006424";
end if;
if first_state_sram_input_id = 6924 then
	sram_write <= x"07DC0020";
end if;
if first_state_sram_input_id = 6925 then
	sram_write <= x"C03C000C";
end if;
if first_state_sram_input_id = 6926 then
	sram_write <= x"C0420008";
end if;
if first_state_sram_input_id = 6927 then
	sram_write <= x"0260FFFF";
end if;
if first_state_sram_input_id = 6928 then
	sram_write <= x"82466CE8";
end if;
if first_state_sram_input_id = 6929 then
	sram_write <= x"22440220";
end if;
if first_state_sram_input_id = 6930 then
	sram_write <= x"C07C0014";
end if;
if first_state_sram_input_id = 6931 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 6932 then
	sram_write <= x"02800000";
end if;
if first_state_sram_input_id = 6933 then
	sram_write <= x"C0BC0000";
end if;
if first_state_sram_input_id = 6934 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 6935 then
	sram_write <= x"006A0000";
end if;
if first_state_sram_input_id = 6936 then
	sram_write <= x"00280000";
end if;
if first_state_sram_input_id = 6937 then
	sram_write <= x"03DC0020";
end if;
if first_state_sram_input_id = 6938 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 6939 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 6940 then
	sram_write <= x"82006424";
end if;
if first_state_sram_input_id = 6941 then
	sram_write <= x"07DC0020";
end if;
if first_state_sram_input_id = 6942 then
	sram_write <= x"C03C000C";
end if;
if first_state_sram_input_id = 6943 then
	sram_write <= x"C042000C";
end if;
if first_state_sram_input_id = 6944 then
	sram_write <= x"0260FFFF";
end if;
if first_state_sram_input_id = 6945 then
	sram_write <= x"82466CE4";
end if;
if first_state_sram_input_id = 6946 then
	sram_write <= x"22440220";
end if;
if first_state_sram_input_id = 6947 then
	sram_write <= x"C07C0014";
end if;
if first_state_sram_input_id = 6948 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 6949 then
	sram_write <= x"02600000";
end if;
if first_state_sram_input_id = 6950 then
	sram_write <= x"C09C0000";
end if;
if first_state_sram_input_id = 6951 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 6952 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 6953 then
	sram_write <= x"00680000";
end if;
if first_state_sram_input_id = 6954 then
	sram_write <= x"03DC0020";
end if;
if first_state_sram_input_id = 6955 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 6956 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 6957 then
	sram_write <= x"82006424";
end if;
if first_state_sram_input_id = 6958 then
	sram_write <= x"07DC0020";
end if;
if first_state_sram_input_id = 6959 then
	sram_write <= x"02200004";
end if;
if first_state_sram_input_id = 6960 then
	sram_write <= x"C05C000C";
end if;
if first_state_sram_input_id = 6961 then
	sram_write <= x"C07C0000";
end if;
if first_state_sram_input_id = 6962 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 6963 then
	sram_write <= x"03DC0020";
end if;
if first_state_sram_input_id = 6964 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 6965 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 6966 then
	sram_write <= x"82006878";
end if;
if first_state_sram_input_id = 6967 then
	sram_write <= x"07DC0020";
end if;
if first_state_sram_input_id = 6968 then
	sram_write <= x"82006CE4";
end if;
if first_state_sram_input_id = 6969 then
	sram_write <= x"82006CE8";
end if;
if first_state_sram_input_id = 6970 then
	sram_write <= x"82006CEC";
end if;
if first_state_sram_input_id = 6971 then
	sram_write <= x"C03C0008";
end if;
if first_state_sram_input_id = 6972 then
	sram_write <= x"02220001";
end if;
if first_state_sram_input_id = 6973 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 6974 then
	sram_write <= x"C07C0004";
end if;
if first_state_sram_input_id = 6975 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 6976 then
	sram_write <= x"C0840000";
end if;
if first_state_sram_input_id = 6977 then
	sram_write <= x"02A0FFFF";
end if;
if first_state_sram_input_id = 6978 then
	sram_write <= x"828A6F84";
end if;
if first_state_sram_input_id = 6979 then
	sram_write <= x"02A00063";
end if;
if first_state_sram_input_id = 6980 then
	sram_write <= x"C43C0018";
end if;
if first_state_sram_input_id = 6981 then
	sram_write <= x"828A6EB4";
end if;
if first_state_sram_input_id = 6982 then
	sram_write <= x"02A000C8";
end if;
if first_state_sram_input_id = 6983 then
	sram_write <= x"22C80220";
end if;
if first_state_sram_input_id = 6984 then
	sram_write <= x"D0AAC000";
end if;
if first_state_sram_input_id = 6985 then
	sram_write <= x"C0CA0028";
end if;
if first_state_sram_input_id = 6986 then
	sram_write <= x"C82C0000";
end if;
if first_state_sram_input_id = 6987 then
	sram_write <= x"C84C0004";
end if;
if first_state_sram_input_id = 6988 then
	sram_write <= x"C86C0008";
end if;
if first_state_sram_input_id = 6989 then
	sram_write <= x"C0FC0000";
end if;
if first_state_sram_input_id = 6990 then
	sram_write <= x"C10E0004";
end if;
if first_state_sram_input_id = 6991 then
	sram_write <= x"22880220";
end if;
if first_state_sram_input_id = 6992 then
	sram_write <= x"D0908000";
end if;
if first_state_sram_input_id = 6993 then
	sram_write <= x"C10A0004";
end if;
if first_state_sram_input_id = 6994 then
	sram_write <= x"03200001";
end if;
if first_state_sram_input_id = 6995 then
	sram_write <= x"C45C001C";
end if;
if first_state_sram_input_id = 6996 then
	sram_write <= x"83126DB0";
end if;
if first_state_sram_input_id = 6997 then
	sram_write <= x"03200002";
end if;
if first_state_sram_input_id = 6998 then
	sram_write <= x"83126D84";
end if;
if first_state_sram_input_id = 6999 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 7000 then
	sram_write <= x"006C0000";
end if;
if first_state_sram_input_id = 7001 then
	sram_write <= x"00480000";
end if;
if first_state_sram_input_id = 7002 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 7003 then
	sram_write <= x"03DC0028";
end if;
if first_state_sram_input_id = 7004 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 7005 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 7006 then
	sram_write <= x"82003BD4";
end if;
if first_state_sram_input_id = 7007 then
	sram_write <= x"07DC0028";
end if;
if first_state_sram_input_id = 7008 then
	sram_write <= x"82006DAC";
end if;
if first_state_sram_input_id = 7009 then
	sram_write <= x"C8280000";
end if;
if first_state_sram_input_id = 7010 then
	sram_write <= x"8E206D94";
end if;
if first_state_sram_input_id = 7011 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 7012 then
	sram_write <= x"82006DAC";
end if;
if first_state_sram_input_id = 7013 then
	sram_write <= x"02A002AC";
end if;
if first_state_sram_input_id = 7014 then
	sram_write <= x"C8280000";
end if;
if first_state_sram_input_id = 7015 then
	sram_write <= x"C84C000C";
end if;
if first_state_sram_input_id = 7016 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 7017 then
	sram_write <= x"CC2A0000";
end if;
if first_state_sram_input_id = 7018 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 7019 then
	sram_write <= x"82006DD8";
end if;
if first_state_sram_input_id = 7020 then
	sram_write <= x"C0CE0000";
end if;
if first_state_sram_input_id = 7021 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 7022 then
	sram_write <= x"00680000";
end if;
if first_state_sram_input_id = 7023 then
	sram_write <= x"004C0000";
end if;
if first_state_sram_input_id = 7024 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 7025 then
	sram_write <= x"03DC0028";
end if;
if first_state_sram_input_id = 7026 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 7027 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 7028 then
	sram_write <= x"8200389C";
end if;
if first_state_sram_input_id = 7029 then
	sram_write <= x"07DC0028";
end if;
if first_state_sram_input_id = 7030 then
	sram_write <= x"82206EB0";
end if;
if first_state_sram_input_id = 7031 then
	sram_write <= x"022002AC";
end if;
if first_state_sram_input_id = 7032 then
	sram_write <= x"C8220000";
end if;
if first_state_sram_input_id = 7033 then
	sram_write <= x"022002B4";
end if;
if first_state_sram_input_id = 7034 then
	sram_write <= x"C8420000";
end if;
if first_state_sram_input_id = 7035 then
	sram_write <= x"8E246DF4";
end if;
if first_state_sram_input_id = 7036 then
	sram_write <= x"82006EAC";
end if;
if first_state_sram_input_id = 7037 then
	sram_write <= x"C03C001C";
end if;
if first_state_sram_input_id = 7038 then
	sram_write <= x"C0420004";
end if;
if first_state_sram_input_id = 7039 then
	sram_write <= x"0260FFFF";
end if;
if first_state_sram_input_id = 7040 then
	sram_write <= x"82466EAC";
end if;
if first_state_sram_input_id = 7041 then
	sram_write <= x"026001E0";
end if;
if first_state_sram_input_id = 7042 then
	sram_write <= x"22440220";
end if;
if first_state_sram_input_id = 7043 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 7044 then
	sram_write <= x"02800000";
end if;
if first_state_sram_input_id = 7045 then
	sram_write <= x"C0BC0000";
end if;
if first_state_sram_input_id = 7046 then
	sram_write <= x"C47C0020";
end if;
if first_state_sram_input_id = 7047 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 7048 then
	sram_write <= x"006A0000";
end if;
if first_state_sram_input_id = 7049 then
	sram_write <= x"00280000";
end if;
if first_state_sram_input_id = 7050 then
	sram_write <= x"03DC002C";
end if;
if first_state_sram_input_id = 7051 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 7052 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 7053 then
	sram_write <= x"82006424";
end if;
if first_state_sram_input_id = 7054 then
	sram_write <= x"07DC002C";
end if;
if first_state_sram_input_id = 7055 then
	sram_write <= x"C03C001C";
end if;
if first_state_sram_input_id = 7056 then
	sram_write <= x"C0420008";
end if;
if first_state_sram_input_id = 7057 then
	sram_write <= x"0260FFFF";
end if;
if first_state_sram_input_id = 7058 then
	sram_write <= x"82466EA8";
end if;
if first_state_sram_input_id = 7059 then
	sram_write <= x"22440220";
end if;
if first_state_sram_input_id = 7060 then
	sram_write <= x"C07C0020";
end if;
if first_state_sram_input_id = 7061 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 7062 then
	sram_write <= x"02600000";
end if;
if first_state_sram_input_id = 7063 then
	sram_write <= x"C09C0000";
end if;
if first_state_sram_input_id = 7064 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 7065 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 7066 then
	sram_write <= x"00680000";
end if;
if first_state_sram_input_id = 7067 then
	sram_write <= x"03DC002C";
end if;
if first_state_sram_input_id = 7068 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 7069 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 7070 then
	sram_write <= x"82006424";
end if;
if first_state_sram_input_id = 7071 then
	sram_write <= x"07DC002C";
end if;
if first_state_sram_input_id = 7072 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 7073 then
	sram_write <= x"C05C001C";
end if;
if first_state_sram_input_id = 7074 then
	sram_write <= x"C07C0000";
end if;
if first_state_sram_input_id = 7075 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 7076 then
	sram_write <= x"03DC002C";
end if;
if first_state_sram_input_id = 7077 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 7078 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 7079 then
	sram_write <= x"82006878";
end if;
if first_state_sram_input_id = 7080 then
	sram_write <= x"07DC002C";
end if;
if first_state_sram_input_id = 7081 then
	sram_write <= x"82006EA8";
end if;
if first_state_sram_input_id = 7082 then
	sram_write <= x"82006EAC";
end if;
if first_state_sram_input_id = 7083 then
	sram_write <= x"82006EB0";
end if;
if first_state_sram_input_id = 7084 then
	sram_write <= x"82006F70";
end if;
if first_state_sram_input_id = 7085 then
	sram_write <= x"C0840004";
end if;
if first_state_sram_input_id = 7086 then
	sram_write <= x"02A0FFFF";
end if;
if first_state_sram_input_id = 7087 then
	sram_write <= x"828A6F70";
end if;
if first_state_sram_input_id = 7088 then
	sram_write <= x"02A001E0";
end if;
if first_state_sram_input_id = 7089 then
	sram_write <= x"22880220";
end if;
if first_state_sram_input_id = 7090 then
	sram_write <= x"D08A8000";
end if;
if first_state_sram_input_id = 7091 then
	sram_write <= x"02C00000";
end if;
if first_state_sram_input_id = 7092 then
	sram_write <= x"C0FC0000";
end if;
if first_state_sram_input_id = 7093 then
	sram_write <= x"C4BC0024";
end if;
if first_state_sram_input_id = 7094 then
	sram_write <= x"C45C001C";
end if;
if first_state_sram_input_id = 7095 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 7096 then
	sram_write <= x"006E0000";
end if;
if first_state_sram_input_id = 7097 then
	sram_write <= x"00480000";
end if;
if first_state_sram_input_id = 7098 then
	sram_write <= x"002C0000";
end if;
if first_state_sram_input_id = 7099 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 7100 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 7101 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 7102 then
	sram_write <= x"82006424";
end if;
if first_state_sram_input_id = 7103 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 7104 then
	sram_write <= x"C03C001C";
end if;
if first_state_sram_input_id = 7105 then
	sram_write <= x"C0420008";
end if;
if first_state_sram_input_id = 7106 then
	sram_write <= x"0260FFFF";
end if;
if first_state_sram_input_id = 7107 then
	sram_write <= x"82466F6C";
end if;
if first_state_sram_input_id = 7108 then
	sram_write <= x"22440220";
end if;
if first_state_sram_input_id = 7109 then
	sram_write <= x"C07C0024";
end if;
if first_state_sram_input_id = 7110 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 7111 then
	sram_write <= x"02600000";
end if;
if first_state_sram_input_id = 7112 then
	sram_write <= x"C09C0000";
end if;
if first_state_sram_input_id = 7113 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 7114 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 7115 then
	sram_write <= x"00680000";
end if;
if first_state_sram_input_id = 7116 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 7117 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 7118 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 7119 then
	sram_write <= x"82006424";
end if;
if first_state_sram_input_id = 7120 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 7121 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 7122 then
	sram_write <= x"C05C001C";
end if;
if first_state_sram_input_id = 7123 then
	sram_write <= x"C07C0000";
end if;
if first_state_sram_input_id = 7124 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 7125 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 7126 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 7127 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 7128 then
	sram_write <= x"82006878";
end if;
if first_state_sram_input_id = 7129 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 7130 then
	sram_write <= x"82006F6C";
end if;
if first_state_sram_input_id = 7131 then
	sram_write <= x"82006F70";
end if;
if first_state_sram_input_id = 7132 then
	sram_write <= x"C03C0018";
end if;
if first_state_sram_input_id = 7133 then
	sram_write <= x"02220001";
end if;
if first_state_sram_input_id = 7134 then
	sram_write <= x"C05C0004";
end if;
if first_state_sram_input_id = 7135 then
	sram_write <= x"C07C0000";
end if;
if first_state_sram_input_id = 7136 then
	sram_write <= x"820069E8";
end if;
if first_state_sram_input_id = 7137 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 7138 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 7139 then
	sram_write <= x"024002B8";
end if;
if first_state_sram_input_id = 7140 then
	sram_write <= x"C8240000";
end if;
if first_state_sram_input_id = 7141 then
	sram_write <= x"C0620014";
end if;
if first_state_sram_input_id = 7142 then
	sram_write <= x"C8460000";
end if;
if first_state_sram_input_id = 7143 then
	sram_write <= x"44224000";
end if;
if first_state_sram_input_id = 7144 then
	sram_write <= x"C8440004";
end if;
if first_state_sram_input_id = 7145 then
	sram_write <= x"C0620014";
end if;
if first_state_sram_input_id = 7146 then
	sram_write <= x"C8660004";
end if;
if first_state_sram_input_id = 7147 then
	sram_write <= x"44446000";
end if;
if first_state_sram_input_id = 7148 then
	sram_write <= x"C8640008";
end if;
if first_state_sram_input_id = 7149 then
	sram_write <= x"C0420014";
end if;
if first_state_sram_input_id = 7150 then
	sram_write <= x"C8840008";
end if;
if first_state_sram_input_id = 7151 then
	sram_write <= x"44668000";
end if;
if first_state_sram_input_id = 7152 then
	sram_write <= x"C0420010";
end if;
if first_state_sram_input_id = 7153 then
	sram_write <= x"C8840000";
end if;
if first_state_sram_input_id = 7154 then
	sram_write <= x"48828000";
end if;
if first_state_sram_input_id = 7155 then
	sram_write <= x"C0420010";
end if;
if first_state_sram_input_id = 7156 then
	sram_write <= x"C8A40004";
end if;
if first_state_sram_input_id = 7157 then
	sram_write <= x"48A4A000";
end if;
if first_state_sram_input_id = 7158 then
	sram_write <= x"C0420010";
end if;
if first_state_sram_input_id = 7159 then
	sram_write <= x"C8C40008";
end if;
if first_state_sram_input_id = 7160 then
	sram_write <= x"48C6C000";
end if;
if first_state_sram_input_id = 7161 then
	sram_write <= x"C042000C";
end if;
if first_state_sram_input_id = 7162 then
	sram_write <= x"C43C0000";
end if;
if first_state_sram_input_id = 7163 then
	sram_write <= x"82407138";
end if;
if first_state_sram_input_id = 7164 then
	sram_write <= x"024002C8";
end if;
if first_state_sram_input_id = 7165 then
	sram_write <= x"C0620024";
end if;
if first_state_sram_input_id = 7166 then
	sram_write <= x"C8E60008";
end if;
if first_state_sram_input_id = 7167 then
	sram_write <= x"48E4E000";
end if;
if first_state_sram_input_id = 7168 then
	sram_write <= x"C0620024";
end if;
if first_state_sram_input_id = 7169 then
	sram_write <= x"C9060004";
end if;
if first_state_sram_input_id = 7170 then
	sram_write <= x"49070000";
end if;
if first_state_sram_input_id = 7171 then
	sram_write <= x"40EF0000";
end if;
if first_state_sram_input_id = 7172 then
	sram_write <= x"C9000080";
end if;
if first_state_sram_input_id = 7173 then
	sram_write <= x"CCDC0008";
end if;
if first_state_sram_input_id = 7174 then
	sram_write <= x"CC5C0010";
end if;
if first_state_sram_input_id = 7175 then
	sram_write <= x"CCBC0018";
end if;
if first_state_sram_input_id = 7176 then
	sram_write <= x"CD1C0020";
end if;
if first_state_sram_input_id = 7177 then
	sram_write <= x"CC7C0028";
end if;
if first_state_sram_input_id = 7178 then
	sram_write <= x"CC3C0030";
end if;
if first_state_sram_input_id = 7179 then
	sram_write <= x"C45C0038";
end if;
if first_state_sram_input_id = 7180 then
	sram_write <= x"CC9C0040";
end if;
if first_state_sram_input_id = 7181 then
	sram_write <= x"CCFC0048";
end if;
if first_state_sram_input_id = 7182 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 7183 then
	sram_write <= x"40210000";
end if;
if first_state_sram_input_id = 7184 then
	sram_write <= x"03DC0058";
end if;
if first_state_sram_input_id = 7185 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 7186 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 7187 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 7188 then
	sram_write <= x"07DC0058";
end if;
if first_state_sram_input_id = 7189 then
	sram_write <= x"C85C0048";
end if;
if first_state_sram_input_id = 7190 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 7191 then
	sram_write <= x"C85C0040";
end if;
if first_state_sram_input_id = 7192 then
	sram_write <= x"40242000";
end if;
if first_state_sram_input_id = 7193 then
	sram_write <= x"C03C0038";
end if;
if first_state_sram_input_id = 7194 then
	sram_write <= x"CC220000";
end if;
if first_state_sram_input_id = 7195 then
	sram_write <= x"C05C0000";
end if;
if first_state_sram_input_id = 7196 then
	sram_write <= x"C0640024";
end if;
if first_state_sram_input_id = 7197 then
	sram_write <= x"C8260008";
end if;
if first_state_sram_input_id = 7198 then
	sram_write <= x"C85C0030";
end if;
if first_state_sram_input_id = 7199 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 7200 then
	sram_write <= x"C0640024";
end if;
if first_state_sram_input_id = 7201 then
	sram_write <= x"C8660000";
end if;
if first_state_sram_input_id = 7202 then
	sram_write <= x"C89C0028";
end if;
if first_state_sram_input_id = 7203 then
	sram_write <= x"48686000";
end if;
if first_state_sram_input_id = 7204 then
	sram_write <= x"40226000";
end if;
if first_state_sram_input_id = 7205 then
	sram_write <= x"C87C0020";
end if;
if first_state_sram_input_id = 7206 then
	sram_write <= x"CC3C0050";
end if;
if first_state_sram_input_id = 7207 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 7208 then
	sram_write <= x"40206000";
end if;
if first_state_sram_input_id = 7209 then
	sram_write <= x"03DC0060";
end if;
if first_state_sram_input_id = 7210 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 7211 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 7212 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 7213 then
	sram_write <= x"07DC0060";
end if;
if first_state_sram_input_id = 7214 then
	sram_write <= x"C85C0050";
end if;
if first_state_sram_input_id = 7215 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 7216 then
	sram_write <= x"C85C0018";
end if;
if first_state_sram_input_id = 7217 then
	sram_write <= x"40242000";
end if;
if first_state_sram_input_id = 7218 then
	sram_write <= x"C03C0038";
end if;
if first_state_sram_input_id = 7219 then
	sram_write <= x"CC220004";
end if;
if first_state_sram_input_id = 7220 then
	sram_write <= x"C05C0000";
end if;
if first_state_sram_input_id = 7221 then
	sram_write <= x"C0640024";
end if;
if first_state_sram_input_id = 7222 then
	sram_write <= x"C8260004";
end if;
if first_state_sram_input_id = 7223 then
	sram_write <= x"C85C0030";
end if;
if first_state_sram_input_id = 7224 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 7225 then
	sram_write <= x"C0640024";
end if;
if first_state_sram_input_id = 7226 then
	sram_write <= x"C8460000";
end if;
if first_state_sram_input_id = 7227 then
	sram_write <= x"C87C0010";
end if;
if first_state_sram_input_id = 7228 then
	sram_write <= x"48464000";
end if;
if first_state_sram_input_id = 7229 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 7230 then
	sram_write <= x"C85C0020";
end if;
if first_state_sram_input_id = 7231 then
	sram_write <= x"CC3C0058";
end if;
if first_state_sram_input_id = 7232 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 7233 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 7234 then
	sram_write <= x"03DC0068";
end if;
if first_state_sram_input_id = 7235 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 7236 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 7237 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 7238 then
	sram_write <= x"07DC0068";
end if;
if first_state_sram_input_id = 7239 then
	sram_write <= x"C85C0058";
end if;
if first_state_sram_input_id = 7240 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 7241 then
	sram_write <= x"C85C0008";
end if;
if first_state_sram_input_id = 7242 then
	sram_write <= x"40242000";
end if;
if first_state_sram_input_id = 7243 then
	sram_write <= x"C03C0038";
end if;
if first_state_sram_input_id = 7244 then
	sram_write <= x"CC220008";
end if;
if first_state_sram_input_id = 7245 then
	sram_write <= x"82007148";
end if;
if first_state_sram_input_id = 7246 then
	sram_write <= x"024002C8";
end if;
if first_state_sram_input_id = 7247 then
	sram_write <= x"CC840000";
end if;
if first_state_sram_input_id = 7248 then
	sram_write <= x"CCA40004";
end if;
if first_state_sram_input_id = 7249 then
	sram_write <= x"CCC40008";
end if;
if first_state_sram_input_id = 7250 then
	sram_write <= x"022002C8";
end if;
if first_state_sram_input_id = 7251 then
	sram_write <= x"C05C0000";
end if;
if first_state_sram_input_id = 7252 then
	sram_write <= x"C0440018";
end if;
if first_state_sram_input_id = 7253 then
	sram_write <= x"8200161C";
end if;
if first_state_sram_input_id = 7254 then
	sram_write <= x"C0620000";
end if;
if first_state_sram_input_id = 7255 then
	sram_write <= x"028002D4";
end if;
if first_state_sram_input_id = 7256 then
	sram_write <= x"C0A20020";
end if;
if first_state_sram_input_id = 7257 then
	sram_write <= x"C82A0000";
end if;
if first_state_sram_input_id = 7258 then
	sram_write <= x"CC280000";
end if;
if first_state_sram_input_id = 7259 then
	sram_write <= x"C0A20020";
end if;
if first_state_sram_input_id = 7260 then
	sram_write <= x"C82A0004";
end if;
if first_state_sram_input_id = 7261 then
	sram_write <= x"CC280004";
end if;
if first_state_sram_input_id = 7262 then
	sram_write <= x"C0A20020";
end if;
if first_state_sram_input_id = 7263 then
	sram_write <= x"C82A0008";
end if;
if first_state_sram_input_id = 7264 then
	sram_write <= x"CC280008";
end if;
if first_state_sram_input_id = 7265 then
	sram_write <= x"02A00001";
end if;
if first_state_sram_input_id = 7266 then
	sram_write <= x"826A7710";
end if;
if first_state_sram_input_id = 7267 then
	sram_write <= x"02A00002";
end if;
if first_state_sram_input_id = 7268 then
	sram_write <= x"826A7648";
end if;
if first_state_sram_input_id = 7269 then
	sram_write <= x"02A00003";
end if;
if first_state_sram_input_id = 7270 then
	sram_write <= x"826A74E8";
end if;
if first_state_sram_input_id = 7271 then
	sram_write <= x"02A00004";
end if;
if first_state_sram_input_id = 7272 then
	sram_write <= x"826A71A8";
end if;
if first_state_sram_input_id = 7273 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 7274 then
	sram_write <= x"C8240000";
end if;
if first_state_sram_input_id = 7275 then
	sram_write <= x"C0620014";
end if;
if first_state_sram_input_id = 7276 then
	sram_write <= x"C8460000";
end if;
if first_state_sram_input_id = 7277 then
	sram_write <= x"44224000";
end if;
if first_state_sram_input_id = 7278 then
	sram_write <= x"C0620010";
end if;
if first_state_sram_input_id = 7279 then
	sram_write <= x"C8460000";
end if;
if first_state_sram_input_id = 7280 then
	sram_write <= x"C49C0000";
end if;
if first_state_sram_input_id = 7281 then
	sram_write <= x"C43C0004";
end if;
if first_state_sram_input_id = 7282 then
	sram_write <= x"C45C0008";
end if;
if first_state_sram_input_id = 7283 then
	sram_write <= x"CC3C0010";
end if;
if first_state_sram_input_id = 7284 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 7285 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 7286 then
	sram_write <= x"03DC0020";
end if;
if first_state_sram_input_id = 7287 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 7288 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 7289 then
	sram_write <= x"8200083C";
end if;
if first_state_sram_input_id = 7290 then
	sram_write <= x"07DC0020";
end if;
if first_state_sram_input_id = 7291 then
	sram_write <= x"C85C0010";
end if;
if first_state_sram_input_id = 7292 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 7293 then
	sram_write <= x"C03C0008";
end if;
if first_state_sram_input_id = 7294 then
	sram_write <= x"C8420008";
end if;
if first_state_sram_input_id = 7295 then
	sram_write <= x"C05C0004";
end if;
if first_state_sram_input_id = 7296 then
	sram_write <= x"C0640014";
end if;
if first_state_sram_input_id = 7297 then
	sram_write <= x"C8660008";
end if;
if first_state_sram_input_id = 7298 then
	sram_write <= x"44446000";
end if;
if first_state_sram_input_id = 7299 then
	sram_write <= x"C0640010";
end if;
if first_state_sram_input_id = 7300 then
	sram_write <= x"C8660008";
end if;
if first_state_sram_input_id = 7301 then
	sram_write <= x"CC3C0018";
end if;
if first_state_sram_input_id = 7302 then
	sram_write <= x"CC5C0020";
end if;
if first_state_sram_input_id = 7303 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 7304 then
	sram_write <= x"40206000";
end if;
if first_state_sram_input_id = 7305 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 7306 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 7307 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 7308 then
	sram_write <= x"8200083C";
end if;
if first_state_sram_input_id = 7309 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 7310 then
	sram_write <= x"C85C0020";
end if;
if first_state_sram_input_id = 7311 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 7312 then
	sram_write <= x"C85C0018";
end if;
if first_state_sram_input_id = 7313 then
	sram_write <= x"48644000";
end if;
if first_state_sram_input_id = 7314 then
	sram_write <= x"48822000";
end if;
if first_state_sram_input_id = 7315 then
	sram_write <= x"40668000";
end if;
if first_state_sram_input_id = 7316 then
	sram_write <= x"8E40725C";
end if;
if first_state_sram_input_id = 7317 then
	sram_write <= x"40804000";
end if;
if first_state_sram_input_id = 7318 then
	sram_write <= x"82007260";
end if;
if first_state_sram_input_id = 7319 then
	sram_write <= x"44804000";
end if;
if first_state_sram_input_id = 7320 then
	sram_write <= x"C8A0006C";
end if;
if first_state_sram_input_id = 7321 then
	sram_write <= x"CCBC0028";
end if;
if first_state_sram_input_id = 7322 then
	sram_write <= x"CC7C0030";
end if;
if first_state_sram_input_id = 7323 then
	sram_write <= x"8E8A7310";
end if;
if first_state_sram_input_id = 7324 then
	sram_write <= x"CC3C0038";
end if;
if first_state_sram_input_id = 7325 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 7326 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 7327 then
	sram_write <= x"03DC0048";
end if;
if first_state_sram_input_id = 7328 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 7329 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 7330 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 7331 then
	sram_write <= x"07DC0048";
end if;
if first_state_sram_input_id = 7332 then
	sram_write <= x"C85C0038";
end if;
if first_state_sram_input_id = 7333 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 7334 then
	sram_write <= x"8E2072A0";
end if;
if first_state_sram_input_id = 7335 then
	sram_write <= x"820072A4";
end if;
if first_state_sram_input_id = 7336 then
	sram_write <= x"44202000";
end if;
if first_state_sram_input_id = 7337 then
	sram_write <= x"C8400068";
end if;
if first_state_sram_input_id = 7338 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 7339 then
	sram_write <= x"C8600064";
end if;
if first_state_sram_input_id = 7340 then
	sram_write <= x"44446000";
end if;
if first_state_sram_input_id = 7341 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 7342 then
	sram_write <= x"C8600060";
end if;
if first_state_sram_input_id = 7343 then
	sram_write <= x"44446000";
end if;
if first_state_sram_input_id = 7344 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 7345 then
	sram_write <= x"C860005C";
end if;
if first_state_sram_input_id = 7346 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 7347 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 7348 then
	sram_write <= x"C8400058";
end if;
if first_state_sram_input_id = 7349 then
	sram_write <= x"44224000";
end if;
if first_state_sram_input_id = 7350 then
	sram_write <= x"C8400054";
end if;
if first_state_sram_input_id = 7351 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 7352 then
	sram_write <= x"C8400050";
end if;
if first_state_sram_input_id = 7353 then
	sram_write <= x"CC3C0040";
end if;
if first_state_sram_input_id = 7354 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 7355 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 7356 then
	sram_write <= x"03DC0050";
end if;
if first_state_sram_input_id = 7357 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 7358 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 7359 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 7360 then
	sram_write <= x"07DC0050";
end if;
if first_state_sram_input_id = 7361 then
	sram_write <= x"C85C0040";
end if;
if first_state_sram_input_id = 7362 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 7363 then
	sram_write <= x"82007314";
end if;
if first_state_sram_input_id = 7364 then
	sram_write <= x"C820004C";
end if;
if first_state_sram_input_id = 7365 then
	sram_write <= x"54220000";
end if;
if first_state_sram_input_id = 7366 then
	sram_write <= x"8E027338";
end if;
if first_state_sram_input_id = 7367 then
	sram_write <= x"58420000";
end if;
if first_state_sram_input_id = 7368 then
	sram_write <= x"8A427330";
end if;
if first_state_sram_input_id = 7369 then
	sram_write <= x"06220001";
end if;
if first_state_sram_input_id = 7370 then
	sram_write <= x"58420000";
end if;
if first_state_sram_input_id = 7371 then
	sram_write <= x"82007334";
end if;
if first_state_sram_input_id = 7372 then
	sram_write <= x"40402000";
end if;
if first_state_sram_input_id = 7373 then
	sram_write <= x"8200733C";
end if;
if first_state_sram_input_id = 7374 then
	sram_write <= x"58420000";
end if;
if first_state_sram_input_id = 7375 then
	sram_write <= x"44224000";
end if;
if first_state_sram_input_id = 7376 then
	sram_write <= x"C03C0008";
end if;
if first_state_sram_input_id = 7377 then
	sram_write <= x"C8420004";
end if;
if first_state_sram_input_id = 7378 then
	sram_write <= x"C03C0004";
end if;
if first_state_sram_input_id = 7379 then
	sram_write <= x"C0420014";
end if;
if first_state_sram_input_id = 7380 then
	sram_write <= x"C8640004";
end if;
if first_state_sram_input_id = 7381 then
	sram_write <= x"44446000";
end if;
if first_state_sram_input_id = 7382 then
	sram_write <= x"C0220010";
end if;
if first_state_sram_input_id = 7383 then
	sram_write <= x"C8620004";
end if;
if first_state_sram_input_id = 7384 then
	sram_write <= x"CC3C0048";
end if;
if first_state_sram_input_id = 7385 then
	sram_write <= x"CC5C0050";
end if;
if first_state_sram_input_id = 7386 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 7387 then
	sram_write <= x"40206000";
end if;
if first_state_sram_input_id = 7388 then
	sram_write <= x"03DC0060";
end if;
if first_state_sram_input_id = 7389 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 7390 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 7391 then
	sram_write <= x"8200083C";
end if;
if first_state_sram_input_id = 7392 then
	sram_write <= x"07DC0060";
end if;
if first_state_sram_input_id = 7393 then
	sram_write <= x"C85C0050";
end if;
if first_state_sram_input_id = 7394 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 7395 then
	sram_write <= x"C85C0030";
end if;
if first_state_sram_input_id = 7396 then
	sram_write <= x"8E40739C";
end if;
if first_state_sram_input_id = 7397 then
	sram_write <= x"40604000";
end if;
if first_state_sram_input_id = 7398 then
	sram_write <= x"820073A0";
end if;
if first_state_sram_input_id = 7399 then
	sram_write <= x"44604000";
end if;
if first_state_sram_input_id = 7400 then
	sram_write <= x"C89C0028";
end if;
if first_state_sram_input_id = 7401 then
	sram_write <= x"8E687448";
end if;
if first_state_sram_input_id = 7402 then
	sram_write <= x"CC3C0058";
end if;
if first_state_sram_input_id = 7403 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 7404 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 7405 then
	sram_write <= x"03DC0068";
end if;
if first_state_sram_input_id = 7406 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 7407 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 7408 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 7409 then
	sram_write <= x"07DC0068";
end if;
if first_state_sram_input_id = 7410 then
	sram_write <= x"C85C0058";
end if;
if first_state_sram_input_id = 7411 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 7412 then
	sram_write <= x"8E2073D8";
end if;
if first_state_sram_input_id = 7413 then
	sram_write <= x"820073DC";
end if;
if first_state_sram_input_id = 7414 then
	sram_write <= x"44202000";
end if;
if first_state_sram_input_id = 7415 then
	sram_write <= x"C8400068";
end if;
if first_state_sram_input_id = 7416 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 7417 then
	sram_write <= x"C8600064";
end if;
if first_state_sram_input_id = 7418 then
	sram_write <= x"44446000";
end if;
if first_state_sram_input_id = 7419 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 7420 then
	sram_write <= x"C8600060";
end if;
if first_state_sram_input_id = 7421 then
	sram_write <= x"44446000";
end if;
if first_state_sram_input_id = 7422 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 7423 then
	sram_write <= x"C860005C";
end if;
if first_state_sram_input_id = 7424 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 7425 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 7426 then
	sram_write <= x"C8400058";
end if;
if first_state_sram_input_id = 7427 then
	sram_write <= x"44224000";
end if;
if first_state_sram_input_id = 7428 then
	sram_write <= x"C8400054";
end if;
if first_state_sram_input_id = 7429 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 7430 then
	sram_write <= x"C8400050";
end if;
if first_state_sram_input_id = 7431 then
	sram_write <= x"CC3C0060";
end if;
if first_state_sram_input_id = 7432 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 7433 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 7434 then
	sram_write <= x"03DC0070";
end if;
if first_state_sram_input_id = 7435 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 7436 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 7437 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 7438 then
	sram_write <= x"07DC0070";
end if;
if first_state_sram_input_id = 7439 then
	sram_write <= x"C85C0060";
end if;
if first_state_sram_input_id = 7440 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 7441 then
	sram_write <= x"8200744C";
end if;
if first_state_sram_input_id = 7442 then
	sram_write <= x"C820004C";
end if;
if first_state_sram_input_id = 7443 then
	sram_write <= x"54220000";
end if;
if first_state_sram_input_id = 7444 then
	sram_write <= x"8E027470";
end if;
if first_state_sram_input_id = 7445 then
	sram_write <= x"58420000";
end if;
if first_state_sram_input_id = 7446 then
	sram_write <= x"8A427468";
end if;
if first_state_sram_input_id = 7447 then
	sram_write <= x"06220001";
end if;
if first_state_sram_input_id = 7448 then
	sram_write <= x"58420000";
end if;
if first_state_sram_input_id = 7449 then
	sram_write <= x"8200746C";
end if;
if first_state_sram_input_id = 7450 then
	sram_write <= x"40402000";
end if;
if first_state_sram_input_id = 7451 then
	sram_write <= x"82007474";
end if;
if first_state_sram_input_id = 7452 then
	sram_write <= x"58420000";
end if;
if first_state_sram_input_id = 7453 then
	sram_write <= x"44224000";
end if;
if first_state_sram_input_id = 7454 then
	sram_write <= x"C8400048";
end if;
if first_state_sram_input_id = 7455 then
	sram_write <= x"C86000A4";
end if;
if first_state_sram_input_id = 7456 then
	sram_write <= x"C89C0048";
end if;
if first_state_sram_input_id = 7457 then
	sram_write <= x"44868000";
end if;
if first_state_sram_input_id = 7458 then
	sram_write <= x"48888000";
end if;
if first_state_sram_input_id = 7459 then
	sram_write <= x"44448000";
end if;
if first_state_sram_input_id = 7460 then
	sram_write <= x"44262000";
end if;
if first_state_sram_input_id = 7461 then
	sram_write <= x"48222000";
end if;
if first_state_sram_input_id = 7462 then
	sram_write <= x"44242000";
end if;
if first_state_sram_input_id = 7463 then
	sram_write <= x"8E2074A4";
end if;
if first_state_sram_input_id = 7464 then
	sram_write <= x"820074A8";
end if;
if first_state_sram_input_id = 7465 then
	sram_write <= x"40200000";
end if;
if first_state_sram_input_id = 7466 then
	sram_write <= x"C8400044";
end if;
if first_state_sram_input_id = 7467 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 7468 then
	sram_write <= x"C8400040";
end if;
if first_state_sram_input_id = 7469 then
	sram_write <= x"CC3C0068";
end if;
if first_state_sram_input_id = 7470 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 7471 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 7472 then
	sram_write <= x"03DC0078";
end if;
if first_state_sram_input_id = 7473 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 7474 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 7475 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 7476 then
	sram_write <= x"07DC0078";
end if;
if first_state_sram_input_id = 7477 then
	sram_write <= x"C85C0068";
end if;
if first_state_sram_input_id = 7478 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 7479 then
	sram_write <= x"C03C0000";
end if;
if first_state_sram_input_id = 7480 then
	sram_write <= x"CC220008";
end if;
if first_state_sram_input_id = 7481 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 7482 then
	sram_write <= x"C8240000";
end if;
if first_state_sram_input_id = 7483 then
	sram_write <= x"C0620014";
end if;
if first_state_sram_input_id = 7484 then
	sram_write <= x"C8460000";
end if;
if first_state_sram_input_id = 7485 then
	sram_write <= x"44224000";
end if;
if first_state_sram_input_id = 7486 then
	sram_write <= x"C8440008";
end if;
if first_state_sram_input_id = 7487 then
	sram_write <= x"C0220014";
end if;
if first_state_sram_input_id = 7488 then
	sram_write <= x"C8620008";
end if;
if first_state_sram_input_id = 7489 then
	sram_write <= x"44446000";
end if;
if first_state_sram_input_id = 7490 then
	sram_write <= x"48222000";
end if;
if first_state_sram_input_id = 7491 then
	sram_write <= x"48444000";
end if;
if first_state_sram_input_id = 7492 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 7493 then
	sram_write <= x"C49C0000";
end if;
if first_state_sram_input_id = 7494 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 7495 then
	sram_write <= x"03DC0078";
end if;
if first_state_sram_input_id = 7496 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 7497 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 7498 then
	sram_write <= x"8200083C";
end if;
if first_state_sram_input_id = 7499 then
	sram_write <= x"07DC0078";
end if;
if first_state_sram_input_id = 7500 then
	sram_write <= x"C840003C";
end if;
if first_state_sram_input_id = 7501 then
	sram_write <= x"CC3C0070";
end if;
if first_state_sram_input_id = 7502 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 7503 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 7504 then
	sram_write <= x"03DC0080";
end if;
if first_state_sram_input_id = 7505 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 7506 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 7507 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 7508 then
	sram_write <= x"07DC0080";
end if;
if first_state_sram_input_id = 7509 then
	sram_write <= x"C85C0070";
end if;
if first_state_sram_input_id = 7510 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 7511 then
	sram_write <= x"54220000";
end if;
if first_state_sram_input_id = 7512 then
	sram_write <= x"8E027580";
end if;
if first_state_sram_input_id = 7513 then
	sram_write <= x"58420000";
end if;
if first_state_sram_input_id = 7514 then
	sram_write <= x"8A427578";
end if;
if first_state_sram_input_id = 7515 then
	sram_write <= x"06220001";
end if;
if first_state_sram_input_id = 7516 then
	sram_write <= x"58420000";
end if;
if first_state_sram_input_id = 7517 then
	sram_write <= x"8200757C";
end if;
if first_state_sram_input_id = 7518 then
	sram_write <= x"40402000";
end if;
if first_state_sram_input_id = 7519 then
	sram_write <= x"82007584";
end if;
if first_state_sram_input_id = 7520 then
	sram_write <= x"58420000";
end if;
if first_state_sram_input_id = 7521 then
	sram_write <= x"44224000";
end if;
if first_state_sram_input_id = 7522 then
	sram_write <= x"C8400050";
end if;
if first_state_sram_input_id = 7523 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 7524 then
	sram_write <= x"C8400098";
end if;
if first_state_sram_input_id = 7525 then
	sram_write <= x"8E2475B8";
end if;
if first_state_sram_input_id = 7526 then
	sram_write <= x"44224000";
end if;
if first_state_sram_input_id = 7527 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 7528 then
	sram_write <= x"03DC0080";
end if;
if first_state_sram_input_id = 7529 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 7530 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 7531 then
	sram_write <= x"82001270";
end if;
if first_state_sram_input_id = 7532 then
	sram_write <= x"07DC0080";
end if;
if first_state_sram_input_id = 7533 then
	sram_write <= x"82007620";
end if;
if first_state_sram_input_id = 7534 then
	sram_write <= x"8E027604";
end if;
if first_state_sram_input_id = 7535 then
	sram_write <= x"C8600090";
end if;
if first_state_sram_input_id = 7536 then
	sram_write <= x"8E6275E4";
end if;
if first_state_sram_input_id = 7537 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 7538 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 7539 then
	sram_write <= x"03DC0080";
end if;
if first_state_sram_input_id = 7540 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 7541 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 7542 then
	sram_write <= x"82001270";
end if;
if first_state_sram_input_id = 7543 then
	sram_write <= x"07DC0080";
end if;
if first_state_sram_input_id = 7544 then
	sram_write <= x"82007600";
end if;
if first_state_sram_input_id = 7545 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 7546 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 7547 then
	sram_write <= x"03DC0080";
end if;
if first_state_sram_input_id = 7548 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 7549 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 7550 then
	sram_write <= x"82000B88";
end if;
if first_state_sram_input_id = 7551 then
	sram_write <= x"07DC0080";
end if;
if first_state_sram_input_id = 7552 then
	sram_write <= x"82007620";
end if;
if first_state_sram_input_id = 7553 then
	sram_write <= x"0220FFFF";
end if;
if first_state_sram_input_id = 7554 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 7555 then
	sram_write <= x"03DC0080";
end if;
if first_state_sram_input_id = 7556 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 7557 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 7558 then
	sram_write <= x"82000B88";
end if;
if first_state_sram_input_id = 7559 then
	sram_write <= x"07DC0080";
end if;
if first_state_sram_input_id = 7560 then
	sram_write <= x"48222000";
end if;
if first_state_sram_input_id = 7561 then
	sram_write <= x"C8400044";
end if;
if first_state_sram_input_id = 7562 then
	sram_write <= x"48624000";
end if;
if first_state_sram_input_id = 7563 then
	sram_write <= x"C03C0000";
end if;
if first_state_sram_input_id = 7564 then
	sram_write <= x"CC620004";
end if;
if first_state_sram_input_id = 7565 then
	sram_write <= x"C86000A8";
end if;
if first_state_sram_input_id = 7566 then
	sram_write <= x"44262000";
end if;
if first_state_sram_input_id = 7567 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 7568 then
	sram_write <= x"CC220008";
end if;
if first_state_sram_input_id = 7569 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 7570 then
	sram_write <= x"C8240004";
end if;
if first_state_sram_input_id = 7571 then
	sram_write <= x"C8400038";
end if;
if first_state_sram_input_id = 7572 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 7573 then
	sram_write <= x"C8400098";
end if;
if first_state_sram_input_id = 7574 then
	sram_write <= x"C49C0000";
end if;
if first_state_sram_input_id = 7575 then
	sram_write <= x"8E247680";
end if;
if first_state_sram_input_id = 7576 then
	sram_write <= x"44224000";
end if;
if first_state_sram_input_id = 7577 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 7578 then
	sram_write <= x"03DC0080";
end if;
if first_state_sram_input_id = 7579 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 7580 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 7581 then
	sram_write <= x"82000EC4";
end if;
if first_state_sram_input_id = 7582 then
	sram_write <= x"07DC0080";
end if;
if first_state_sram_input_id = 7583 then
	sram_write <= x"820076E8";
end if;
if first_state_sram_input_id = 7584 then
	sram_write <= x"8E0276CC";
end if;
if first_state_sram_input_id = 7585 then
	sram_write <= x"C8600090";
end if;
if first_state_sram_input_id = 7586 then
	sram_write <= x"8E6276AC";
end if;
if first_state_sram_input_id = 7587 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 7588 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 7589 then
	sram_write <= x"03DC0080";
end if;
if first_state_sram_input_id = 7590 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 7591 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 7592 then
	sram_write <= x"82000EC4";
end if;
if first_state_sram_input_id = 7593 then
	sram_write <= x"07DC0080";
end if;
if first_state_sram_input_id = 7594 then
	sram_write <= x"820076C8";
end if;
if first_state_sram_input_id = 7595 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 7596 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 7597 then
	sram_write <= x"03DC0080";
end if;
if first_state_sram_input_id = 7598 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 7599 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 7600 then
	sram_write <= x"8200084C";
end if;
if first_state_sram_input_id = 7601 then
	sram_write <= x"07DC0080";
end if;
if first_state_sram_input_id = 7602 then
	sram_write <= x"820076E8";
end if;
if first_state_sram_input_id = 7603 then
	sram_write <= x"0220FFFF";
end if;
if first_state_sram_input_id = 7604 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 7605 then
	sram_write <= x"03DC0080";
end if;
if first_state_sram_input_id = 7606 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 7607 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 7608 then
	sram_write <= x"8200084C";
end if;
if first_state_sram_input_id = 7609 then
	sram_write <= x"07DC0080";
end if;
if first_state_sram_input_id = 7610 then
	sram_write <= x"48222000";
end if;
if first_state_sram_input_id = 7611 then
	sram_write <= x"C8400044";
end if;
if first_state_sram_input_id = 7612 then
	sram_write <= x"48642000";
end if;
if first_state_sram_input_id = 7613 then
	sram_write <= x"C03C0000";
end if;
if first_state_sram_input_id = 7614 then
	sram_write <= x"CC620000";
end if;
if first_state_sram_input_id = 7615 then
	sram_write <= x"C86000A8";
end if;
if first_state_sram_input_id = 7616 then
	sram_write <= x"44262000";
end if;
if first_state_sram_input_id = 7617 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 7618 then
	sram_write <= x"CC220004";
end if;
if first_state_sram_input_id = 7619 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 7620 then
	sram_write <= x"C8240000";
end if;
if first_state_sram_input_id = 7621 then
	sram_write <= x"C0620014";
end if;
if first_state_sram_input_id = 7622 then
	sram_write <= x"C8460000";
end if;
if first_state_sram_input_id = 7623 then
	sram_write <= x"44224000";
end if;
if first_state_sram_input_id = 7624 then
	sram_write <= x"C8400034";
end if;
if first_state_sram_input_id = 7625 then
	sram_write <= x"48624000";
end if;
if first_state_sram_input_id = 7626 then
	sram_write <= x"54660000";
end if;
if first_state_sram_input_id = 7627 then
	sram_write <= x"8E067748";
end if;
if first_state_sram_input_id = 7628 then
	sram_write <= x"58860000";
end if;
if first_state_sram_input_id = 7629 then
	sram_write <= x"8A867744";
end if;
if first_state_sram_input_id = 7630 then
	sram_write <= x"06660001";
end if;
if first_state_sram_input_id = 7631 then
	sram_write <= x"58660000";
end if;
if first_state_sram_input_id = 7632 then
	sram_write <= x"82007744";
end if;
if first_state_sram_input_id = 7633 then
	sram_write <= x"8200774C";
end if;
if first_state_sram_input_id = 7634 then
	sram_write <= x"58660000";
end if;
if first_state_sram_input_id = 7635 then
	sram_write <= x"C8800030";
end if;
if first_state_sram_input_id = 7636 then
	sram_write <= x"48668000";
end if;
if first_state_sram_input_id = 7637 then
	sram_write <= x"44226000";
end if;
if first_state_sram_input_id = 7638 then
	sram_write <= x"C860003C";
end if;
if first_state_sram_input_id = 7639 then
	sram_write <= x"C8A40008";
end if;
if first_state_sram_input_id = 7640 then
	sram_write <= x"C0220014";
end if;
if first_state_sram_input_id = 7641 then
	sram_write <= x"C8C20008";
end if;
if first_state_sram_input_id = 7642 then
	sram_write <= x"44AAC000";
end if;
if first_state_sram_input_id = 7643 then
	sram_write <= x"484A4000";
end if;
if first_state_sram_input_id = 7644 then
	sram_write <= x"54240000";
end if;
if first_state_sram_input_id = 7645 then
	sram_write <= x"8E047790";
end if;
if first_state_sram_input_id = 7646 then
	sram_write <= x"58C20000";
end if;
if first_state_sram_input_id = 7647 then
	sram_write <= x"8AC4778C";
end if;
if first_state_sram_input_id = 7648 then
	sram_write <= x"06220001";
end if;
if first_state_sram_input_id = 7649 then
	sram_write <= x"58420000";
end if;
if first_state_sram_input_id = 7650 then
	sram_write <= x"8200778C";
end if;
if first_state_sram_input_id = 7651 then
	sram_write <= x"82007794";
end if;
if first_state_sram_input_id = 7652 then
	sram_write <= x"58420000";
end if;
if first_state_sram_input_id = 7653 then
	sram_write <= x"48448000";
end if;
if first_state_sram_input_id = 7654 then
	sram_write <= x"444A4000";
end if;
if first_state_sram_input_id = 7655 then
	sram_write <= x"8E2677B4";
end if;
if first_state_sram_input_id = 7656 then
	sram_write <= x"8E4677AC";
end if;
if first_state_sram_input_id = 7657 then
	sram_write <= x"C8200044";
end if;
if first_state_sram_input_id = 7658 then
	sram_write <= x"820077B0";
end if;
if first_state_sram_input_id = 7659 then
	sram_write <= x"40200000";
end if;
if first_state_sram_input_id = 7660 then
	sram_write <= x"820077C4";
end if;
if first_state_sram_input_id = 7661 then
	sram_write <= x"8E4677C0";
end if;
if first_state_sram_input_id = 7662 then
	sram_write <= x"40200000";
end if;
if first_state_sram_input_id = 7663 then
	sram_write <= x"820077C4";
end if;
if first_state_sram_input_id = 7664 then
	sram_write <= x"C8200044";
end if;
if first_state_sram_input_id = 7665 then
	sram_write <= x"CC280004";
end if;
if first_state_sram_input_id = 7666 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 7667 then
	sram_write <= x"8E0277D4";
end if;
if first_state_sram_input_id = 7668 then
	sram_write <= x"82007818";
end if;
if first_state_sram_input_id = 7669 then
	sram_write <= x"022002EC";
end if;
if first_state_sram_input_id = 7670 then
	sram_write <= x"024002D4";
end if;
if first_state_sram_input_id = 7671 then
	sram_write <= x"C8820000";
end if;
if first_state_sram_input_id = 7672 then
	sram_write <= x"C8A40000";
end if;
if first_state_sram_input_id = 7673 then
	sram_write <= x"48A2A000";
end if;
if first_state_sram_input_id = 7674 then
	sram_write <= x"4088A000";
end if;
if first_state_sram_input_id = 7675 then
	sram_write <= x"CC820000";
end if;
if first_state_sram_input_id = 7676 then
	sram_write <= x"C8820004";
end if;
if first_state_sram_input_id = 7677 then
	sram_write <= x"C8A40004";
end if;
if first_state_sram_input_id = 7678 then
	sram_write <= x"48A2A000";
end if;
if first_state_sram_input_id = 7679 then
	sram_write <= x"4088A000";
end if;
if first_state_sram_input_id = 7680 then
	sram_write <= x"CC820004";
end if;
if first_state_sram_input_id = 7681 then
	sram_write <= x"C8820008";
end if;
if first_state_sram_input_id = 7682 then
	sram_write <= x"C8A40008";
end if;
if first_state_sram_input_id = 7683 then
	sram_write <= x"4822A000";
end if;
if first_state_sram_input_id = 7684 then
	sram_write <= x"40282000";
end if;
if first_state_sram_input_id = 7685 then
	sram_write <= x"CC220008";
end if;
if first_state_sram_input_id = 7686 then
	sram_write <= x"8E047820";
end if;
if first_state_sram_input_id = 7687 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 7688 then
	sram_write <= x"48244000";
end if;
if first_state_sram_input_id = 7689 then
	sram_write <= x"48222000";
end if;
if first_state_sram_input_id = 7690 then
	sram_write <= x"48226000";
end if;
if first_state_sram_input_id = 7691 then
	sram_write <= x"022002EC";
end if;
if first_state_sram_input_id = 7692 then
	sram_write <= x"C8420000";
end if;
if first_state_sram_input_id = 7693 then
	sram_write <= x"40442000";
end if;
if first_state_sram_input_id = 7694 then
	sram_write <= x"CC420000";
end if;
if first_state_sram_input_id = 7695 then
	sram_write <= x"C8420004";
end if;
if first_state_sram_input_id = 7696 then
	sram_write <= x"40442000";
end if;
if first_state_sram_input_id = 7697 then
	sram_write <= x"CC420004";
end if;
if first_state_sram_input_id = 7698 then
	sram_write <= x"C8420008";
end if;
if first_state_sram_input_id = 7699 then
	sram_write <= x"40242000";
end if;
if first_state_sram_input_id = 7700 then
	sram_write <= x"CC220008";
end if;
if first_state_sram_input_id = 7701 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 7702 then
	sram_write <= x"86207A10";
end if;
if first_state_sram_input_id = 7703 then
	sram_write <= x"02600370";
end if;
if first_state_sram_input_id = 7704 then
	sram_write <= x"22820220";
end if;
if first_state_sram_input_id = 7705 then
	sram_write <= x"D0668000";
end if;
if first_state_sram_input_id = 7706 then
	sram_write <= x"C0860004";
end if;
if first_state_sram_input_id = 7707 then
	sram_write <= x"02A002B4";
end if;
if first_state_sram_input_id = 7708 then
	sram_write <= x"C860002C";
end if;
if first_state_sram_input_id = 7709 then
	sram_write <= x"CC6A0000";
end if;
if first_state_sram_input_id = 7710 then
	sram_write <= x"02C00000";
end if;
if first_state_sram_input_id = 7711 then
	sram_write <= x"02E002A8";
end if;
if first_state_sram_input_id = 7712 then
	sram_write <= x"C10E0000";
end if;
if first_state_sram_input_id = 7713 then
	sram_write <= x"C43C0000";
end if;
if first_state_sram_input_id = 7714 then
	sram_write <= x"CC5C0008";
end if;
if first_state_sram_input_id = 7715 then
	sram_write <= x"C45C0010";
end if;
if first_state_sram_input_id = 7716 then
	sram_write <= x"CC3C0018";
end if;
if first_state_sram_input_id = 7717 then
	sram_write <= x"C49C0020";
end if;
if first_state_sram_input_id = 7718 then
	sram_write <= x"C4FC0024";
end if;
if first_state_sram_input_id = 7719 then
	sram_write <= x"C47C0028";
end if;
if first_state_sram_input_id = 7720 then
	sram_write <= x"C4BC002C";
end if;
if first_state_sram_input_id = 7721 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 7722 then
	sram_write <= x"00680000";
end if;
if first_state_sram_input_id = 7723 then
	sram_write <= x"00500000";
end if;
if first_state_sram_input_id = 7724 then
	sram_write <= x"002C0000";
end if;
if first_state_sram_input_id = 7725 then
	sram_write <= x"03DC0038";
end if;
if first_state_sram_input_id = 7726 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 7727 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 7728 then
	sram_write <= x"820069E8";
end if;
if first_state_sram_input_id = 7729 then
	sram_write <= x"07DC0038";
end if;
if first_state_sram_input_id = 7730 then
	sram_write <= x"C03C002C";
end if;
if first_state_sram_input_id = 7731 then
	sram_write <= x"C8220000";
end if;
if first_state_sram_input_id = 7732 then
	sram_write <= x"C8400070";
end if;
if first_state_sram_input_id = 7733 then
	sram_write <= x"8E4278E0";
end if;
if first_state_sram_input_id = 7734 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 7735 then
	sram_write <= x"820078F4";
end if;
if first_state_sram_input_id = 7736 then
	sram_write <= x"C8400028";
end if;
if first_state_sram_input_id = 7737 then
	sram_write <= x"8E2478F0";
end if;
if first_state_sram_input_id = 7738 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 7739 then
	sram_write <= x"820078F4";
end if;
if first_state_sram_input_id = 7740 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 7741 then
	sram_write <= x"822079F8";
end if;
if first_state_sram_input_id = 7742 then
	sram_write <= x"022002C4";
end if;
if first_state_sram_input_id = 7743 then
	sram_write <= x"C0220000";
end if;
if first_state_sram_input_id = 7744 then
	sram_write <= x"22220220";
end if;
if first_state_sram_input_id = 7745 then
	sram_write <= x"024002B0";
end if;
if first_state_sram_input_id = 7746 then
	sram_write <= x"C0440000";
end if;
if first_state_sram_input_id = 7747 then
	sram_write <= x"00224000";
end if;
if first_state_sram_input_id = 7748 then
	sram_write <= x"C05C0028";
end if;
if first_state_sram_input_id = 7749 then
	sram_write <= x"C0640000";
end if;
if first_state_sram_input_id = 7750 then
	sram_write <= x"82267920";
end if;
if first_state_sram_input_id = 7751 then
	sram_write <= x"820079F4";
end if;
if first_state_sram_input_id = 7752 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 7753 then
	sram_write <= x"C07C0024";
end if;
if first_state_sram_input_id = 7754 then
	sram_write <= x"C0660000";
end if;
if first_state_sram_input_id = 7755 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 7756 then
	sram_write <= x"00460000";
end if;
if first_state_sram_input_id = 7757 then
	sram_write <= x"03DC0038";
end if;
if first_state_sram_input_id = 7758 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 7759 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 7760 then
	sram_write <= x"82005414";
end if;
if first_state_sram_input_id = 7761 then
	sram_write <= x"07DC0038";
end if;
if first_state_sram_input_id = 7762 then
	sram_write <= x"82207950";
end if;
if first_state_sram_input_id = 7763 then
	sram_write <= x"820079F4";
end if;
if first_state_sram_input_id = 7764 then
	sram_write <= x"022002C8";
end if;
if first_state_sram_input_id = 7765 then
	sram_write <= x"C05C0020";
end if;
if first_state_sram_input_id = 7766 then
	sram_write <= x"C0640000";
end if;
if first_state_sram_input_id = 7767 then
	sram_write <= x"C8220000";
end if;
if first_state_sram_input_id = 7768 then
	sram_write <= x"C8460000";
end if;
if first_state_sram_input_id = 7769 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 7770 then
	sram_write <= x"C8420004";
end if;
if first_state_sram_input_id = 7771 then
	sram_write <= x"C8660004";
end if;
if first_state_sram_input_id = 7772 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 7773 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 7774 then
	sram_write <= x"C8420008";
end if;
if first_state_sram_input_id = 7775 then
	sram_write <= x"C8660008";
end if;
if first_state_sram_input_id = 7776 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 7777 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 7778 then
	sram_write <= x"C03C0028";
end if;
if first_state_sram_input_id = 7779 then
	sram_write <= x"C8420008";
end if;
if first_state_sram_input_id = 7780 then
	sram_write <= x"C87C0018";
end if;
if first_state_sram_input_id = 7781 then
	sram_write <= x"48846000";
end if;
if first_state_sram_input_id = 7782 then
	sram_write <= x"48282000";
end if;
if first_state_sram_input_id = 7783 then
	sram_write <= x"C0240000";
end if;
if first_state_sram_input_id = 7784 then
	sram_write <= x"C05C0010";
end if;
if first_state_sram_input_id = 7785 then
	sram_write <= x"C8840000";
end if;
if first_state_sram_input_id = 7786 then
	sram_write <= x"C8A20000";
end if;
if first_state_sram_input_id = 7787 then
	sram_write <= x"4888A000";
end if;
if first_state_sram_input_id = 7788 then
	sram_write <= x"C8A40004";
end if;
if first_state_sram_input_id = 7789 then
	sram_write <= x"C8C20004";
end if;
if first_state_sram_input_id = 7790 then
	sram_write <= x"48AAC000";
end if;
if first_state_sram_input_id = 7791 then
	sram_write <= x"4088A000";
end if;
if first_state_sram_input_id = 7792 then
	sram_write <= x"C8A40008";
end if;
if first_state_sram_input_id = 7793 then
	sram_write <= x"C8C20008";
end if;
if first_state_sram_input_id = 7794 then
	sram_write <= x"48AAC000";
end if;
if first_state_sram_input_id = 7795 then
	sram_write <= x"4088A000";
end if;
if first_state_sram_input_id = 7796 then
	sram_write <= x"48448000";
end if;
if first_state_sram_input_id = 7797 then
	sram_write <= x"C89C0008";
end if;
if first_state_sram_input_id = 7798 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 7799 then
	sram_write <= x"40608000";
end if;
if first_state_sram_input_id = 7800 then
	sram_write <= x"03DC0038";
end if;
if first_state_sram_input_id = 7801 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 7802 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 7803 then
	sram_write <= x"820077CC";
end if;
if first_state_sram_input_id = 7804 then
	sram_write <= x"07DC0038";
end if;
if first_state_sram_input_id = 7805 then
	sram_write <= x"820079F8";
end if;
if first_state_sram_input_id = 7806 then
	sram_write <= x"C03C0000";
end if;
if first_state_sram_input_id = 7807 then
	sram_write <= x"06220001";
end if;
if first_state_sram_input_id = 7808 then
	sram_write <= x"C83C0018";
end if;
if first_state_sram_input_id = 7809 then
	sram_write <= x"C85C0008";
end if;
if first_state_sram_input_id = 7810 then
	sram_write <= x"C05C0010";
end if;
if first_state_sram_input_id = 7811 then
	sram_write <= x"82007858";
end if;
if first_state_sram_input_id = 7812 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 7813 then
	sram_write <= x"02800004";
end if;
if first_state_sram_input_id = 7814 then
	sram_write <= x"86828030";
end if;
if first_state_sram_input_id = 7815 then
	sram_write <= x"C0860008";
end if;
if first_state_sram_input_id = 7816 then
	sram_write <= x"02A002B4";
end if;
if first_state_sram_input_id = 7817 then
	sram_write <= x"C860002C";
end if;
if first_state_sram_input_id = 7818 then
	sram_write <= x"CC6A0000";
end if;
if first_state_sram_input_id = 7819 then
	sram_write <= x"02C00000";
end if;
if first_state_sram_input_id = 7820 then
	sram_write <= x"02E002A8";
end if;
if first_state_sram_input_id = 7821 then
	sram_write <= x"C10E0000";
end if;
if first_state_sram_input_id = 7822 then
	sram_write <= x"CC5C0000";
end if;
if first_state_sram_input_id = 7823 then
	sram_write <= x"C4FC0008";
end if;
if first_state_sram_input_id = 7824 then
	sram_write <= x"C47C000C";
end if;
if first_state_sram_input_id = 7825 then
	sram_write <= x"CC3C0010";
end if;
if first_state_sram_input_id = 7826 then
	sram_write <= x"C45C0018";
end if;
if first_state_sram_input_id = 7827 then
	sram_write <= x"C49C001C";
end if;
if first_state_sram_input_id = 7828 then
	sram_write <= x"C43C0020";
end if;
if first_state_sram_input_id = 7829 then
	sram_write <= x"C4BC0024";
end if;
if first_state_sram_input_id = 7830 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 7831 then
	sram_write <= x"00640000";
end if;
if first_state_sram_input_id = 7832 then
	sram_write <= x"002C0000";
end if;
if first_state_sram_input_id = 7833 then
	sram_write <= x"00500000";
end if;
if first_state_sram_input_id = 7834 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 7835 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 7836 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 7837 then
	sram_write <= x"82005E4C";
end if;
if first_state_sram_input_id = 7838 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 7839 then
	sram_write <= x"C03C0024";
end if;
if first_state_sram_input_id = 7840 then
	sram_write <= x"C8220000";
end if;
if first_state_sram_input_id = 7841 then
	sram_write <= x"C8400070";
end if;
if first_state_sram_input_id = 7842 then
	sram_write <= x"8E427A94";
end if;
if first_state_sram_input_id = 7843 then
	sram_write <= x"02400000";
end if;
if first_state_sram_input_id = 7844 then
	sram_write <= x"82007AA8";
end if;
if first_state_sram_input_id = 7845 then
	sram_write <= x"C8400028";
end if;
if first_state_sram_input_id = 7846 then
	sram_write <= x"8E247AA4";
end if;
if first_state_sram_input_id = 7847 then
	sram_write <= x"02400000";
end if;
if first_state_sram_input_id = 7848 then
	sram_write <= x"82007AA8";
end if;
if first_state_sram_input_id = 7849 then
	sram_write <= x"02400001";
end if;
if first_state_sram_input_id = 7850 then
	sram_write <= x"82407F8C";
end if;
if first_state_sram_input_id = 7851 then
	sram_write <= x"024002C4";
end if;
if first_state_sram_input_id = 7852 then
	sram_write <= x"C0440000";
end if;
if first_state_sram_input_id = 7853 then
	sram_write <= x"026000C8";
end if;
if first_state_sram_input_id = 7854 then
	sram_write <= x"22840220";
end if;
if first_state_sram_input_id = 7855 then
	sram_write <= x"D0668000";
end if;
if first_state_sram_input_id = 7856 then
	sram_write <= x"C0860008";
end if;
if first_state_sram_input_id = 7857 then
	sram_write <= x"C0A6001C";
end if;
if first_state_sram_input_id = 7858 then
	sram_write <= x"C82A0000";
end if;
if first_state_sram_input_id = 7859 then
	sram_write <= x"C85C0010";
end if;
if first_state_sram_input_id = 7860 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 7861 then
	sram_write <= x"C0A60004";
end if;
if first_state_sram_input_id = 7862 then
	sram_write <= x"02C00001";
end if;
if first_state_sram_input_id = 7863 then
	sram_write <= x"C49C0028";
end if;
if first_state_sram_input_id = 7864 then
	sram_write <= x"CC3C0030";
end if;
if first_state_sram_input_id = 7865 then
	sram_write <= x"C45C0038";
end if;
if first_state_sram_input_id = 7866 then
	sram_write <= x"C47C003C";
end if;
if first_state_sram_input_id = 7867 then
	sram_write <= x"82AC7B50";
end if;
if first_state_sram_input_id = 7868 then
	sram_write <= x"02C00002";
end if;
if first_state_sram_input_id = 7869 then
	sram_write <= x"82AC7B18";
end if;
if first_state_sram_input_id = 7870 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 7871 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 7872 then
	sram_write <= x"03DC0048";
end if;
if first_state_sram_input_id = 7873 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 7874 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 7875 then
	sram_write <= x"82006F8C";
end if;
if first_state_sram_input_id = 7876 then
	sram_write <= x"07DC0048";
end if;
if first_state_sram_input_id = 7877 then
	sram_write <= x"82007B4C";
end if;
if first_state_sram_input_id = 7878 then
	sram_write <= x"02A002C8";
end if;
if first_state_sram_input_id = 7879 then
	sram_write <= x"C0C60010";
end if;
if first_state_sram_input_id = 7880 then
	sram_write <= x"C86C0000";
end if;
if first_state_sram_input_id = 7881 then
	sram_write <= x"44606000";
end if;
if first_state_sram_input_id = 7882 then
	sram_write <= x"CC6A0000";
end if;
if first_state_sram_input_id = 7883 then
	sram_write <= x"C0C60010";
end if;
if first_state_sram_input_id = 7884 then
	sram_write <= x"C86C0004";
end if;
if first_state_sram_input_id = 7885 then
	sram_write <= x"44606000";
end if;
if first_state_sram_input_id = 7886 then
	sram_write <= x"CC6A0004";
end if;
if first_state_sram_input_id = 7887 then
	sram_write <= x"C0C60010";
end if;
if first_state_sram_input_id = 7888 then
	sram_write <= x"C86C0008";
end if;
if first_state_sram_input_id = 7889 then
	sram_write <= x"44606000";
end if;
if first_state_sram_input_id = 7890 then
	sram_write <= x"CC6A0008";
end if;
if first_state_sram_input_id = 7891 then
	sram_write <= x"82007BA4";
end if;
if first_state_sram_input_id = 7892 then
	sram_write <= x"02A002B0";
end if;
if first_state_sram_input_id = 7893 then
	sram_write <= x"C0AA0000";
end if;
if first_state_sram_input_id = 7894 then
	sram_write <= x"02C002C8";
end if;
if first_state_sram_input_id = 7895 then
	sram_write <= x"CC0C0000";
end if;
if first_state_sram_input_id = 7896 then
	sram_write <= x"CC0C0004";
end if;
if first_state_sram_input_id = 7897 then
	sram_write <= x"CC0C0008";
end if;
if first_state_sram_input_id = 7898 then
	sram_write <= x"06EA0001";
end if;
if first_state_sram_input_id = 7899 then
	sram_write <= x"06AA0001";
end if;
if first_state_sram_input_id = 7900 then
	sram_write <= x"22AA0220";
end if;
if first_state_sram_input_id = 7901 then
	sram_write <= x"C11C0018";
end if;
if first_state_sram_input_id = 7902 then
	sram_write <= x"D870A000";
end if;
if first_state_sram_input_id = 7903 then
	sram_write <= x"8A607B94";
end if;
if first_state_sram_input_id = 7904 then
	sram_write <= x"8E067B8C";
end if;
if first_state_sram_input_id = 7905 then
	sram_write <= x"C860007C";
end if;
if first_state_sram_input_id = 7906 then
	sram_write <= x"82007B90";
end if;
if first_state_sram_input_id = 7907 then
	sram_write <= x"C86000A8";
end if;
if first_state_sram_input_id = 7908 then
	sram_write <= x"82007B98";
end if;
if first_state_sram_input_id = 7909 then
	sram_write <= x"40600000";
end if;
if first_state_sram_input_id = 7910 then
	sram_write <= x"44606000";
end if;
if first_state_sram_input_id = 7911 then
	sram_write <= x"22AE0220";
end if;
if first_state_sram_input_id = 7912 then
	sram_write <= x"DC6CA000";
end if;
if first_state_sram_input_id = 7913 then
	sram_write <= x"0220030C";
end if;
if first_state_sram_input_id = 7914 then
	sram_write <= x"024002B8";
end if;
if first_state_sram_input_id = 7915 then
	sram_write <= x"C8240000";
end if;
if first_state_sram_input_id = 7916 then
	sram_write <= x"CC220000";
end if;
if first_state_sram_input_id = 7917 then
	sram_write <= x"C8240004";
end if;
if first_state_sram_input_id = 7918 then
	sram_write <= x"CC220004";
end if;
if first_state_sram_input_id = 7919 then
	sram_write <= x"C8240008";
end if;
if first_state_sram_input_id = 7920 then
	sram_write <= x"CC220008";
end if;
if first_state_sram_input_id = 7921 then
	sram_write <= x"C03C003C";
end if;
if first_state_sram_input_id = 7922 then
	sram_write <= x"C45C0040";
end if;
if first_state_sram_input_id = 7923 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 7924 then
	sram_write <= x"03DC004C";
end if;
if first_state_sram_input_id = 7925 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 7926 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 7927 then
	sram_write <= x"82007158";
end if;
if first_state_sram_input_id = 7928 then
	sram_write <= x"07DC004C";
end if;
if first_state_sram_input_id = 7929 then
	sram_write <= x"C03C0038";
end if;
if first_state_sram_input_id = 7930 then
	sram_write <= x"22220220";
end if;
if first_state_sram_input_id = 7931 then
	sram_write <= x"024002B0";
end if;
if first_state_sram_input_id = 7932 then
	sram_write <= x"C0440000";
end if;
if first_state_sram_input_id = 7933 then
	sram_write <= x"00224000";
end if;
if first_state_sram_input_id = 7934 then
	sram_write <= x"C05C0020";
end if;
if first_state_sram_input_id = 7935 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 7936 then
	sram_write <= x"C09C001C";
end if;
if first_state_sram_input_id = 7937 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 7938 then
	sram_write <= x"C03C000C";
end if;
if first_state_sram_input_id = 7939 then
	sram_write <= x"C0620004";
end if;
if first_state_sram_input_id = 7940 then
	sram_write <= x"22A40220";
end if;
if first_state_sram_input_id = 7941 then
	sram_write <= x"D066A000";
end if;
if first_state_sram_input_id = 7942 then
	sram_write <= x"C0BC0040";
end if;
if first_state_sram_input_id = 7943 then
	sram_write <= x"C82A0000";
end if;
if first_state_sram_input_id = 7944 then
	sram_write <= x"CC260000";
end if;
if first_state_sram_input_id = 7945 then
	sram_write <= x"C82A0004";
end if;
if first_state_sram_input_id = 7946 then
	sram_write <= x"CC260004";
end if;
if first_state_sram_input_id = 7947 then
	sram_write <= x"C82A0008";
end if;
if first_state_sram_input_id = 7948 then
	sram_write <= x"CC260008";
end if;
if first_state_sram_input_id = 7949 then
	sram_write <= x"C062000C";
end if;
if first_state_sram_input_id = 7950 then
	sram_write <= x"C0DC003C";
end if;
if first_state_sram_input_id = 7951 then
	sram_write <= x"C0EC001C";
end if;
if first_state_sram_input_id = 7952 then
	sram_write <= x"C82E0000";
end if;
if first_state_sram_input_id = 7953 then
	sram_write <= x"C84000A4";
end if;
if first_state_sram_input_id = 7954 then
	sram_write <= x"8E247D0C";
end if;
if first_state_sram_input_id = 7955 then
	sram_write <= x"02E00001";
end if;
if first_state_sram_input_id = 7956 then
	sram_write <= x"23040220";
end if;
if first_state_sram_input_id = 7957 then
	sram_write <= x"D4E70000";
end if;
if first_state_sram_input_id = 7958 then
	sram_write <= x"C0620010";
end if;
if first_state_sram_input_id = 7959 then
	sram_write <= x"22E40220";
end if;
if first_state_sram_input_id = 7960 then
	sram_write <= x"D0E6E000";
end if;
if first_state_sram_input_id = 7961 then
	sram_write <= x"030002D4";
end if;
if first_state_sram_input_id = 7962 then
	sram_write <= x"C8300000";
end if;
if first_state_sram_input_id = 7963 then
	sram_write <= x"CC2E0000";
end if;
if first_state_sram_input_id = 7964 then
	sram_write <= x"C8300004";
end if;
if first_state_sram_input_id = 7965 then
	sram_write <= x"CC2E0004";
end if;
if first_state_sram_input_id = 7966 then
	sram_write <= x"C8300008";
end if;
if first_state_sram_input_id = 7967 then
	sram_write <= x"CC2E0008";
end if;
if first_state_sram_input_id = 7968 then
	sram_write <= x"22E40220";
end if;
if first_state_sram_input_id = 7969 then
	sram_write <= x"D066E000";
end if;
if first_state_sram_input_id = 7970 then
	sram_write <= x"C8200024";
end if;
if first_state_sram_input_id = 7971 then
	sram_write <= x"C47C0044";
end if;
if first_state_sram_input_id = 7972 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 7973 then
	sram_write <= x"03DC0050";
end if;
if first_state_sram_input_id = 7974 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 7975 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 7976 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 7977 then
	sram_write <= x"07DC0050";
end if;
if first_state_sram_input_id = 7978 then
	sram_write <= x"C85C0030";
end if;
if first_state_sram_input_id = 7979 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 7980 then
	sram_write <= x"C03C0044";
end if;
if first_state_sram_input_id = 7981 then
	sram_write <= x"C8620000";
end if;
if first_state_sram_input_id = 7982 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 7983 then
	sram_write <= x"CC620000";
end if;
if first_state_sram_input_id = 7984 then
	sram_write <= x"C8620004";
end if;
if first_state_sram_input_id = 7985 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 7986 then
	sram_write <= x"CC620004";
end if;
if first_state_sram_input_id = 7987 then
	sram_write <= x"C8620008";
end if;
if first_state_sram_input_id = 7988 then
	sram_write <= x"48262000";
end if;
if first_state_sram_input_id = 7989 then
	sram_write <= x"CC220008";
end if;
if first_state_sram_input_id = 7990 then
	sram_write <= x"C03C000C";
end if;
if first_state_sram_input_id = 7991 then
	sram_write <= x"C042001C";
end if;
if first_state_sram_input_id = 7992 then
	sram_write <= x"C07C0020";
end if;
if first_state_sram_input_id = 7993 then
	sram_write <= x"22860220";
end if;
if first_state_sram_input_id = 7994 then
	sram_write <= x"D0448000";
end if;
if first_state_sram_input_id = 7995 then
	sram_write <= x"028002C8";
end if;
if first_state_sram_input_id = 7996 then
	sram_write <= x"C8280000";
end if;
if first_state_sram_input_id = 7997 then
	sram_write <= x"CC240000";
end if;
if first_state_sram_input_id = 7998 then
	sram_write <= x"C8280004";
end if;
if first_state_sram_input_id = 7999 then
	sram_write <= x"CC240004";
end if;
if first_state_sram_input_id = 8000 then
	sram_write <= x"C8280008";
end if;
if first_state_sram_input_id = 8001 then
	sram_write <= x"CC240008";
end if;
if first_state_sram_input_id = 8002 then
	sram_write <= x"82007D18";
end if;
if first_state_sram_input_id = 8003 then
	sram_write <= x"02E00000";
end if;
if first_state_sram_input_id = 8004 then
	sram_write <= x"23040220";
end if;
if first_state_sram_input_id = 8005 then
	sram_write <= x"D4E70000";
end if;
if first_state_sram_input_id = 8006 then
	sram_write <= x"C8200020";
end if;
if first_state_sram_input_id = 8007 then
	sram_write <= x"024002C8";
end if;
if first_state_sram_input_id = 8008 then
	sram_write <= x"C07C0018";
end if;
if first_state_sram_input_id = 8009 then
	sram_write <= x"C8460000";
end if;
if first_state_sram_input_id = 8010 then
	sram_write <= x"C8640000";
end if;
if first_state_sram_input_id = 8011 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 8012 then
	sram_write <= x"C8660004";
end if;
if first_state_sram_input_id = 8013 then
	sram_write <= x"C8840004";
end if;
if first_state_sram_input_id = 8014 then
	sram_write <= x"48668000";
end if;
if first_state_sram_input_id = 8015 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 8016 then
	sram_write <= x"C8660008";
end if;
if first_state_sram_input_id = 8017 then
	sram_write <= x"C8840008";
end if;
if first_state_sram_input_id = 8018 then
	sram_write <= x"48668000";
end if;
if first_state_sram_input_id = 8019 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 8020 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 8021 then
	sram_write <= x"C8460000";
end if;
if first_state_sram_input_id = 8022 then
	sram_write <= x"C8640000";
end if;
if first_state_sram_input_id = 8023 then
	sram_write <= x"48626000";
end if;
if first_state_sram_input_id = 8024 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 8025 then
	sram_write <= x"CC460000";
end if;
if first_state_sram_input_id = 8026 then
	sram_write <= x"C8460004";
end if;
if first_state_sram_input_id = 8027 then
	sram_write <= x"C8640004";
end if;
if first_state_sram_input_id = 8028 then
	sram_write <= x"48626000";
end if;
if first_state_sram_input_id = 8029 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 8030 then
	sram_write <= x"CC460004";
end if;
if first_state_sram_input_id = 8031 then
	sram_write <= x"C8460008";
end if;
if first_state_sram_input_id = 8032 then
	sram_write <= x"C8640008";
end if;
if first_state_sram_input_id = 8033 then
	sram_write <= x"48226000";
end if;
if first_state_sram_input_id = 8034 then
	sram_write <= x"40242000";
end if;
if first_state_sram_input_id = 8035 then
	sram_write <= x"CC260008";
end if;
if first_state_sram_input_id = 8036 then
	sram_write <= x"C09C003C";
end if;
if first_state_sram_input_id = 8037 then
	sram_write <= x"C0A8001C";
end if;
if first_state_sram_input_id = 8038 then
	sram_write <= x"C82A0004";
end if;
if first_state_sram_input_id = 8039 then
	sram_write <= x"C85C0010";
end if;
if first_state_sram_input_id = 8040 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 8041 then
	sram_write <= x"02A00000";
end if;
if first_state_sram_input_id = 8042 then
	sram_write <= x"C0DC0008";
end if;
if first_state_sram_input_id = 8043 then
	sram_write <= x"C0CC0000";
end if;
if first_state_sram_input_id = 8044 then
	sram_write <= x"CC3C0048";
end if;
if first_state_sram_input_id = 8045 then
	sram_write <= x"C45C0050";
end if;
if first_state_sram_input_id = 8046 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 8047 then
	sram_write <= x"004C0000";
end if;
if first_state_sram_input_id = 8048 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 8049 then
	sram_write <= x"03DC005C";
end if;
if first_state_sram_input_id = 8050 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 8051 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 8052 then
	sram_write <= x"82005414";
end if;
if first_state_sram_input_id = 8053 then
	sram_write <= x"07DC005C";
end if;
if first_state_sram_input_id = 8054 then
	sram_write <= x"82207DE0";
end if;
if first_state_sram_input_id = 8055 then
	sram_write <= x"82007E78";
end if;
if first_state_sram_input_id = 8056 then
	sram_write <= x"022001D0";
end if;
if first_state_sram_input_id = 8057 then
	sram_write <= x"C05C0050";
end if;
if first_state_sram_input_id = 8058 then
	sram_write <= x"C8240000";
end if;
if first_state_sram_input_id = 8059 then
	sram_write <= x"C8420000";
end if;
if first_state_sram_input_id = 8060 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 8061 then
	sram_write <= x"C8440004";
end if;
if first_state_sram_input_id = 8062 then
	sram_write <= x"C8620004";
end if;
if first_state_sram_input_id = 8063 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 8064 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 8065 then
	sram_write <= x"C8440008";
end if;
if first_state_sram_input_id = 8066 then
	sram_write <= x"C8620008";
end if;
if first_state_sram_input_id = 8067 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 8068 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 8069 then
	sram_write <= x"44202000";
end if;
if first_state_sram_input_id = 8070 then
	sram_write <= x"C85C0030";
end if;
if first_state_sram_input_id = 8071 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 8072 then
	sram_write <= x"C05C0018";
end if;
if first_state_sram_input_id = 8073 then
	sram_write <= x"C8640000";
end if;
if first_state_sram_input_id = 8074 then
	sram_write <= x"C8820000";
end if;
if first_state_sram_input_id = 8075 then
	sram_write <= x"48668000";
end if;
if first_state_sram_input_id = 8076 then
	sram_write <= x"C8840004";
end if;
if first_state_sram_input_id = 8077 then
	sram_write <= x"C8A20004";
end if;
if first_state_sram_input_id = 8078 then
	sram_write <= x"4888A000";
end if;
if first_state_sram_input_id = 8079 then
	sram_write <= x"40668000";
end if;
if first_state_sram_input_id = 8080 then
	sram_write <= x"C8840008";
end if;
if first_state_sram_input_id = 8081 then
	sram_write <= x"C8A20008";
end if;
if first_state_sram_input_id = 8082 then
	sram_write <= x"4888A000";
end if;
if first_state_sram_input_id = 8083 then
	sram_write <= x"40668000";
end if;
if first_state_sram_input_id = 8084 then
	sram_write <= x"44606000";
end if;
if first_state_sram_input_id = 8085 then
	sram_write <= x"C89C0048";
end if;
if first_state_sram_input_id = 8086 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 8087 then
	sram_write <= x"40406000";
end if;
if first_state_sram_input_id = 8088 then
	sram_write <= x"40608000";
end if;
if first_state_sram_input_id = 8089 then
	sram_write <= x"03DC005C";
end if;
if first_state_sram_input_id = 8090 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 8091 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 8092 then
	sram_write <= x"820077CC";
end if;
if first_state_sram_input_id = 8093 then
	sram_write <= x"07DC005C";
end if;
if first_state_sram_input_id = 8094 then
	sram_write <= x"02200318";
end if;
if first_state_sram_input_id = 8095 then
	sram_write <= x"C05C0040";
end if;
if first_state_sram_input_id = 8096 then
	sram_write <= x"C8240000";
end if;
if first_state_sram_input_id = 8097 then
	sram_write <= x"CC220000";
end if;
if first_state_sram_input_id = 8098 then
	sram_write <= x"C8240004";
end if;
if first_state_sram_input_id = 8099 then
	sram_write <= x"CC220004";
end if;
if first_state_sram_input_id = 8100 then
	sram_write <= x"C8240008";
end if;
if first_state_sram_input_id = 8101 then
	sram_write <= x"CC220008";
end if;
if first_state_sram_input_id = 8102 then
	sram_write <= x"022000C4";
end if;
if first_state_sram_input_id = 8103 then
	sram_write <= x"C0220000";
end if;
if first_state_sram_input_id = 8104 then
	sram_write <= x"06220001";
end if;
if first_state_sram_input_id = 8105 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 8106 then
	sram_write <= x"01240000";
end if;
if first_state_sram_input_id = 8107 then
	sram_write <= x"00420000";
end if;
if first_state_sram_input_id = 8108 then
	sram_write <= x"00320000";
end if;
if first_state_sram_input_id = 8109 then
	sram_write <= x"03DC005C";
end if;
if first_state_sram_input_id = 8110 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 8111 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 8112 then
	sram_write <= x"8200462C";
end if;
if first_state_sram_input_id = 8113 then
	sram_write <= x"07DC005C";
end if;
if first_state_sram_input_id = 8114 then
	sram_write <= x"02200640";
end if;
if first_state_sram_input_id = 8115 then
	sram_write <= x"C0220000";
end if;
if first_state_sram_input_id = 8116 then
	sram_write <= x"06220001";
end if;
if first_state_sram_input_id = 8117 then
	sram_write <= x"C83C0030";
end if;
if first_state_sram_input_id = 8118 then
	sram_write <= x"C85C0048";
end if;
if first_state_sram_input_id = 8119 then
	sram_write <= x"C05C0018";
end if;
if first_state_sram_input_id = 8120 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 8121 then
	sram_write <= x"03DC005C";
end if;
if first_state_sram_input_id = 8122 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 8123 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 8124 then
	sram_write <= x"82007858";
end if;
if first_state_sram_input_id = 8125 then
	sram_write <= x"07DC005C";
end if;
if first_state_sram_input_id = 8126 then
	sram_write <= x"C820001C";
end if;
if first_state_sram_input_id = 8127 then
	sram_write <= x"C85C0010";
end if;
if first_state_sram_input_id = 8128 then
	sram_write <= x"8E247F08";
end if;
if first_state_sram_input_id = 8129 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 8130 then
	sram_write <= x"02200004";
end if;
if first_state_sram_input_id = 8131 then
	sram_write <= x"C05C0020";
end if;
if first_state_sram_input_id = 8132 then
	sram_write <= x"86427F18";
end if;
if first_state_sram_input_id = 8133 then
	sram_write <= x"82007F2C";
end if;
if first_state_sram_input_id = 8134 then
	sram_write <= x"02240001";
end if;
if first_state_sram_input_id = 8135 then
	sram_write <= x"0260FFFF";
end if;
if first_state_sram_input_id = 8136 then
	sram_write <= x"22220220";
end if;
if first_state_sram_input_id = 8137 then
	sram_write <= x"C09C001C";
end if;
if first_state_sram_input_id = 8138 then
	sram_write <= x"D4682000";
end if;
if first_state_sram_input_id = 8139 then
	sram_write <= x"02200002";
end if;
if first_state_sram_input_id = 8140 then
	sram_write <= x"C07C0028";
end if;
if first_state_sram_input_id = 8141 then
	sram_write <= x"82627F3C";
end if;
if first_state_sram_input_id = 8142 then
	sram_write <= x"82007F88";
end if;
if first_state_sram_input_id = 8143 then
	sram_write <= x"C82000A8";
end if;
if first_state_sram_input_id = 8144 then
	sram_write <= x"C03C003C";
end if;
if first_state_sram_input_id = 8145 then
	sram_write <= x"C022001C";
end if;
if first_state_sram_input_id = 8146 then
	sram_write <= x"C8620000";
end if;
if first_state_sram_input_id = 8147 then
	sram_write <= x"44226000";
end if;
if first_state_sram_input_id = 8148 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 8149 then
	sram_write <= x"02240001";
end if;
if first_state_sram_input_id = 8150 then
	sram_write <= x"C05C0024";
end if;
if first_state_sram_input_id = 8151 then
	sram_write <= x"C8440000";
end if;
if first_state_sram_input_id = 8152 then
	sram_write <= x"C87C0000";
end if;
if first_state_sram_input_id = 8153 then
	sram_write <= x"40464000";
end if;
if first_state_sram_input_id = 8154 then
	sram_write <= x"C05C0018";
end if;
if first_state_sram_input_id = 8155 then
	sram_write <= x"C07C000C";
end if;
if first_state_sram_input_id = 8156 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 8157 then
	sram_write <= x"03DC005C";
end if;
if first_state_sram_input_id = 8158 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 8159 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 8160 then
	sram_write <= x"82007A14";
end if;
if first_state_sram_input_id = 8161 then
	sram_write <= x"07DC005C";
end if;
if first_state_sram_input_id = 8162 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 8163 then
	sram_write <= x"0220FFFF";
end if;
if first_state_sram_input_id = 8164 then
	sram_write <= x"C05C0020";
end if;
if first_state_sram_input_id = 8165 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 8166 then
	sram_write <= x"C09C001C";
end if;
if first_state_sram_input_id = 8167 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 8168 then
	sram_write <= x"8240802C";
end if;
if first_state_sram_input_id = 8169 then
	sram_write <= x"022001D0";
end if;
if first_state_sram_input_id = 8170 then
	sram_write <= x"C05C0018";
end if;
if first_state_sram_input_id = 8171 then
	sram_write <= x"C8240000";
end if;
if first_state_sram_input_id = 8172 then
	sram_write <= x"C8420000";
end if;
if first_state_sram_input_id = 8173 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 8174 then
	sram_write <= x"C8440004";
end if;
if first_state_sram_input_id = 8175 then
	sram_write <= x"C8620004";
end if;
if first_state_sram_input_id = 8176 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 8177 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 8178 then
	sram_write <= x"C8440008";
end if;
if first_state_sram_input_id = 8179 then
	sram_write <= x"C8620008";
end if;
if first_state_sram_input_id = 8180 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 8181 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 8182 then
	sram_write <= x"44202000";
end if;
if first_state_sram_input_id = 8183 then
	sram_write <= x"8E027FE4";
end if;
if first_state_sram_input_id = 8184 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 8185 then
	sram_write <= x"48422000";
end if;
if first_state_sram_input_id = 8186 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 8187 then
	sram_write <= x"C85C0010";
end if;
if first_state_sram_input_id = 8188 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 8189 then
	sram_write <= x"022001DC";
end if;
if first_state_sram_input_id = 8190 then
	sram_write <= x"C8420000";
end if;
if first_state_sram_input_id = 8191 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 8192 then
	sram_write <= x"022002EC";
end if;
if first_state_sram_input_id = 8193 then
	sram_write <= x"C8420000";
end if;
if first_state_sram_input_id = 8194 then
	sram_write <= x"40442000";
end if;
if first_state_sram_input_id = 8195 then
	sram_write <= x"CC420000";
end if;
if first_state_sram_input_id = 8196 then
	sram_write <= x"C8420004";
end if;
if first_state_sram_input_id = 8197 then
	sram_write <= x"40442000";
end if;
if first_state_sram_input_id = 8198 then
	sram_write <= x"CC420004";
end if;
if first_state_sram_input_id = 8199 then
	sram_write <= x"C8420008";
end if;
if first_state_sram_input_id = 8200 then
	sram_write <= x"40242000";
end if;
if first_state_sram_input_id = 8201 then
	sram_write <= x"CC220008";
end if;
if first_state_sram_input_id = 8202 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 8203 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 8204 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 8205 then
	sram_write <= x"024002B4";
end if;
if first_state_sram_input_id = 8206 then
	sram_write <= x"C840002C";
end if;
if first_state_sram_input_id = 8207 then
	sram_write <= x"CC440000";
end if;
if first_state_sram_input_id = 8208 then
	sram_write <= x"02600000";
end if;
if first_state_sram_input_id = 8209 then
	sram_write <= x"028002A8";
end if;
if first_state_sram_input_id = 8210 then
	sram_write <= x"C0A80000";
end if;
if first_state_sram_input_id = 8211 then
	sram_write <= x"CC3C0000";
end if;
if first_state_sram_input_id = 8212 then
	sram_write <= x"C49C0008";
end if;
if first_state_sram_input_id = 8213 then
	sram_write <= x"C43C000C";
end if;
if first_state_sram_input_id = 8214 then
	sram_write <= x"C45C0010";
end if;
if first_state_sram_input_id = 8215 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 8216 then
	sram_write <= x"004A0000";
end if;
if first_state_sram_input_id = 8217 then
	sram_write <= x"01260000";
end if;
if first_state_sram_input_id = 8218 then
	sram_write <= x"00620000";
end if;
if first_state_sram_input_id = 8219 then
	sram_write <= x"00320000";
end if;
if first_state_sram_input_id = 8220 then
	sram_write <= x"03DC001C";
end if;
if first_state_sram_input_id = 8221 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 8222 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 8223 then
	sram_write <= x"820069E8";
end if;
if first_state_sram_input_id = 8224 then
	sram_write <= x"07DC001C";
end if;
if first_state_sram_input_id = 8225 then
	sram_write <= x"C03C0010";
end if;
if first_state_sram_input_id = 8226 then
	sram_write <= x"C8220000";
end if;
if first_state_sram_input_id = 8227 then
	sram_write <= x"C8400070";
end if;
if first_state_sram_input_id = 8228 then
	sram_write <= x"8E42809C";
end if;
if first_state_sram_input_id = 8229 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 8230 then
	sram_write <= x"820080B0";
end if;
if first_state_sram_input_id = 8231 then
	sram_write <= x"C8400028";
end if;
if first_state_sram_input_id = 8232 then
	sram_write <= x"8E2480AC";
end if;
if first_state_sram_input_id = 8233 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 8234 then
	sram_write <= x"820080B0";
end if;
if first_state_sram_input_id = 8235 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 8236 then
	sram_write <= x"8220827C";
end if;
if first_state_sram_input_id = 8237 then
	sram_write <= x"022000C8";
end if;
if first_state_sram_input_id = 8238 then
	sram_write <= x"024002C4";
end if;
if first_state_sram_input_id = 8239 then
	sram_write <= x"C0440000";
end if;
if first_state_sram_input_id = 8240 then
	sram_write <= x"22440220";
end if;
if first_state_sram_input_id = 8241 then
	sram_write <= x"D0224000";
end if;
if first_state_sram_input_id = 8242 then
	sram_write <= x"C05C000C";
end if;
if first_state_sram_input_id = 8243 then
	sram_write <= x"C0440000";
end if;
if first_state_sram_input_id = 8244 then
	sram_write <= x"C0620004";
end if;
if first_state_sram_input_id = 8245 then
	sram_write <= x"02800001";
end if;
if first_state_sram_input_id = 8246 then
	sram_write <= x"C43C0014";
end if;
if first_state_sram_input_id = 8247 then
	sram_write <= x"8268813C";
end if;
if first_state_sram_input_id = 8248 then
	sram_write <= x"02400002";
end if;
if first_state_sram_input_id = 8249 then
	sram_write <= x"82648104";
end if;
if first_state_sram_input_id = 8250 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 8251 then
	sram_write <= x"03DC0020";
end if;
if first_state_sram_input_id = 8252 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 8253 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 8254 then
	sram_write <= x"82006F8C";
end if;
if first_state_sram_input_id = 8255 then
	sram_write <= x"07DC0020";
end if;
if first_state_sram_input_id = 8256 then
	sram_write <= x"82008138";
end if;
if first_state_sram_input_id = 8257 then
	sram_write <= x"024002C8";
end if;
if first_state_sram_input_id = 8258 then
	sram_write <= x"C0620010";
end if;
if first_state_sram_input_id = 8259 then
	sram_write <= x"C8260000";
end if;
if first_state_sram_input_id = 8260 then
	sram_write <= x"44202000";
end if;
if first_state_sram_input_id = 8261 then
	sram_write <= x"CC240000";
end if;
if first_state_sram_input_id = 8262 then
	sram_write <= x"C0620010";
end if;
if first_state_sram_input_id = 8263 then
	sram_write <= x"C8260004";
end if;
if first_state_sram_input_id = 8264 then
	sram_write <= x"44202000";
end if;
if first_state_sram_input_id = 8265 then
	sram_write <= x"CC240004";
end if;
if first_state_sram_input_id = 8266 then
	sram_write <= x"C0620010";
end if;
if first_state_sram_input_id = 8267 then
	sram_write <= x"C8260008";
end if;
if first_state_sram_input_id = 8268 then
	sram_write <= x"44202000";
end if;
if first_state_sram_input_id = 8269 then
	sram_write <= x"CC240008";
end if;
if first_state_sram_input_id = 8270 then
	sram_write <= x"8200818C";
end if;
if first_state_sram_input_id = 8271 then
	sram_write <= x"026002B0";
end if;
if first_state_sram_input_id = 8272 then
	sram_write <= x"C0660000";
end if;
if first_state_sram_input_id = 8273 then
	sram_write <= x"028002C8";
end if;
if first_state_sram_input_id = 8274 then
	sram_write <= x"CC080000";
end if;
if first_state_sram_input_id = 8275 then
	sram_write <= x"CC080004";
end if;
if first_state_sram_input_id = 8276 then
	sram_write <= x"CC080008";
end if;
if first_state_sram_input_id = 8277 then
	sram_write <= x"06A60001";
end if;
if first_state_sram_input_id = 8278 then
	sram_write <= x"06660001";
end if;
if first_state_sram_input_id = 8279 then
	sram_write <= x"22660220";
end if;
if first_state_sram_input_id = 8280 then
	sram_write <= x"D8246000";
end if;
if first_state_sram_input_id = 8281 then
	sram_write <= x"8A20817C";
end if;
if first_state_sram_input_id = 8282 then
	sram_write <= x"8E028174";
end if;
if first_state_sram_input_id = 8283 then
	sram_write <= x"C820007C";
end if;
if first_state_sram_input_id = 8284 then
	sram_write <= x"82008178";
end if;
if first_state_sram_input_id = 8285 then
	sram_write <= x"C82000A8";
end if;
if first_state_sram_input_id = 8286 then
	sram_write <= x"82008180";
end if;
if first_state_sram_input_id = 8287 then
	sram_write <= x"40200000";
end if;
if first_state_sram_input_id = 8288 then
	sram_write <= x"44202000";
end if;
if first_state_sram_input_id = 8289 then
	sram_write <= x"224A0220";
end if;
if first_state_sram_input_id = 8290 then
	sram_write <= x"DC284000";
end if;
if first_state_sram_input_id = 8291 then
	sram_write <= x"024002B8";
end if;
if first_state_sram_input_id = 8292 then
	sram_write <= x"C03C0014";
end if;
if first_state_sram_input_id = 8293 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 8294 then
	sram_write <= x"03DC0020";
end if;
if first_state_sram_input_id = 8295 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 8296 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 8297 then
	sram_write <= x"82007158";
end if;
if first_state_sram_input_id = 8298 then
	sram_write <= x"07DC0020";
end if;
if first_state_sram_input_id = 8299 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 8300 then
	sram_write <= x"C05C0008";
end if;
if first_state_sram_input_id = 8301 then
	sram_write <= x"C0440000";
end if;
if first_state_sram_input_id = 8302 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 8303 then
	sram_write <= x"03DC0020";
end if;
if first_state_sram_input_id = 8304 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 8305 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 8306 then
	sram_write <= x"82005414";
end if;
if first_state_sram_input_id = 8307 then
	sram_write <= x"07DC0020";
end if;
if first_state_sram_input_id = 8308 then
	sram_write <= x"822081D8";
end if;
if first_state_sram_input_id = 8309 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 8310 then
	sram_write <= x"022002C8";
end if;
if first_state_sram_input_id = 8311 then
	sram_write <= x"024001D0";
end if;
if first_state_sram_input_id = 8312 then
	sram_write <= x"C8220000";
end if;
if first_state_sram_input_id = 8313 then
	sram_write <= x"C8440000";
end if;
if first_state_sram_input_id = 8314 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 8315 then
	sram_write <= x"C8420004";
end if;
if first_state_sram_input_id = 8316 then
	sram_write <= x"C8640004";
end if;
if first_state_sram_input_id = 8317 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 8318 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 8319 then
	sram_write <= x"C8420008";
end if;
if first_state_sram_input_id = 8320 then
	sram_write <= x"C8640008";
end if;
if first_state_sram_input_id = 8321 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 8322 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 8323 then
	sram_write <= x"44202000";
end if;
if first_state_sram_input_id = 8324 then
	sram_write <= x"8E02821C";
end if;
if first_state_sram_input_id = 8325 then
	sram_write <= x"40200000";
end if;
if first_state_sram_input_id = 8326 then
	sram_write <= x"8200821C";
end if;
if first_state_sram_input_id = 8327 then
	sram_write <= x"022002E0";
end if;
if first_state_sram_input_id = 8328 then
	sram_write <= x"C85C0000";
end if;
if first_state_sram_input_id = 8329 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 8330 then
	sram_write <= x"C05C0014";
end if;
if first_state_sram_input_id = 8331 then
	sram_write <= x"C044001C";
end if;
if first_state_sram_input_id = 8332 then
	sram_write <= x"C8440000";
end if;
if first_state_sram_input_id = 8333 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 8334 then
	sram_write <= x"024002D4";
end if;
if first_state_sram_input_id = 8335 then
	sram_write <= x"C8420000";
end if;
if first_state_sram_input_id = 8336 then
	sram_write <= x"C8640000";
end if;
if first_state_sram_input_id = 8337 then
	sram_write <= x"48626000";
end if;
if first_state_sram_input_id = 8338 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 8339 then
	sram_write <= x"CC420000";
end if;
if first_state_sram_input_id = 8340 then
	sram_write <= x"C8420004";
end if;
if first_state_sram_input_id = 8341 then
	sram_write <= x"C8640004";
end if;
if first_state_sram_input_id = 8342 then
	sram_write <= x"48626000";
end if;
if first_state_sram_input_id = 8343 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 8344 then
	sram_write <= x"CC420004";
end if;
if first_state_sram_input_id = 8345 then
	sram_write <= x"C8420008";
end if;
if first_state_sram_input_id = 8346 then
	sram_write <= x"C8640008";
end if;
if first_state_sram_input_id = 8347 then
	sram_write <= x"48226000";
end if;
if first_state_sram_input_id = 8348 then
	sram_write <= x"40242000";
end if;
if first_state_sram_input_id = 8349 then
	sram_write <= x"CC220008";
end if;
if first_state_sram_input_id = 8350 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 8351 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 8352 then
	sram_write <= x"86808490";
end if;
if first_state_sram_input_id = 8353 then
	sram_write <= x"22A80220";
end if;
if first_state_sram_input_id = 8354 then
	sram_write <= x"D0A2A000";
end if;
if first_state_sram_input_id = 8355 then
	sram_write <= x"C0CA0000";
end if;
if first_state_sram_input_id = 8356 then
	sram_write <= x"C82C0000";
end if;
if first_state_sram_input_id = 8357 then
	sram_write <= x"C8440000";
end if;
if first_state_sram_input_id = 8358 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 8359 then
	sram_write <= x"C84C0004";
end if;
if first_state_sram_input_id = 8360 then
	sram_write <= x"C8640004";
end if;
if first_state_sram_input_id = 8361 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 8362 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 8363 then
	sram_write <= x"C84C0008";
end if;
if first_state_sram_input_id = 8364 then
	sram_write <= x"C8640008";
end if;
if first_state_sram_input_id = 8365 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 8366 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 8367 then
	sram_write <= x"C47C0000";
end if;
if first_state_sram_input_id = 8368 then
	sram_write <= x"C45C0004";
end if;
if first_state_sram_input_id = 8369 then
	sram_write <= x"C43C0008";
end if;
if first_state_sram_input_id = 8370 then
	sram_write <= x"C49C000C";
end if;
if first_state_sram_input_id = 8371 then
	sram_write <= x"8E208320";
end if;
if first_state_sram_input_id = 8372 then
	sram_write <= x"C8400018";
end if;
if first_state_sram_input_id = 8373 then
	sram_write <= x"C4BC0010";
end if;
if first_state_sram_input_id = 8374 then
	sram_write <= x"CC3C0018";
end if;
if first_state_sram_input_id = 8375 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 8376 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 8377 then
	sram_write <= x"03DC0028";
end if;
if first_state_sram_input_id = 8378 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 8379 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 8380 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 8381 then
	sram_write <= x"07DC0028";
end if;
if first_state_sram_input_id = 8382 then
	sram_write <= x"C85C0018";
end if;
if first_state_sram_input_id = 8383 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 8384 then
	sram_write <= x"C03C0010";
end if;
if first_state_sram_input_id = 8385 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 8386 then
	sram_write <= x"03DC0028";
end if;
if first_state_sram_input_id = 8387 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 8388 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 8389 then
	sram_write <= x"82008034";
end if;
if first_state_sram_input_id = 8390 then
	sram_write <= x"07DC0028";
end if;
if first_state_sram_input_id = 8391 then
	sram_write <= x"82008378";
end if;
if first_state_sram_input_id = 8392 then
	sram_write <= x"02A80001";
end if;
if first_state_sram_input_id = 8393 then
	sram_write <= x"22AA0220";
end if;
if first_state_sram_input_id = 8394 then
	sram_write <= x"D0A2A000";
end if;
if first_state_sram_input_id = 8395 then
	sram_write <= x"C8400014";
end if;
if first_state_sram_input_id = 8396 then
	sram_write <= x"C4BC0020";
end if;
if first_state_sram_input_id = 8397 then
	sram_write <= x"CC3C0018";
end if;
if first_state_sram_input_id = 8398 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 8399 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 8400 then
	sram_write <= x"03DC002C";
end if;
if first_state_sram_input_id = 8401 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 8402 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 8403 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 8404 then
	sram_write <= x"07DC002C";
end if;
if first_state_sram_input_id = 8405 then
	sram_write <= x"C85C0018";
end if;
if first_state_sram_input_id = 8406 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 8407 then
	sram_write <= x"C03C0020";
end if;
if first_state_sram_input_id = 8408 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 8409 then
	sram_write <= x"03DC002C";
end if;
if first_state_sram_input_id = 8410 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 8411 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 8412 then
	sram_write <= x"82008034";
end if;
if first_state_sram_input_id = 8413 then
	sram_write <= x"07DC002C";
end if;
if first_state_sram_input_id = 8414 then
	sram_write <= x"C03C000C";
end if;
if first_state_sram_input_id = 8415 then
	sram_write <= x"06220002";
end if;
if first_state_sram_input_id = 8416 then
	sram_write <= x"8620848C";
end if;
if first_state_sram_input_id = 8417 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 8418 then
	sram_write <= x"C07C0008";
end if;
if first_state_sram_input_id = 8419 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 8420 then
	sram_write <= x"C0840000";
end if;
if first_state_sram_input_id = 8421 then
	sram_write <= x"C8280000";
end if;
if first_state_sram_input_id = 8422 then
	sram_write <= x"C0BC0004";
end if;
if first_state_sram_input_id = 8423 then
	sram_write <= x"C84A0000";
end if;
if first_state_sram_input_id = 8424 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 8425 then
	sram_write <= x"C8480004";
end if;
if first_state_sram_input_id = 8426 then
	sram_write <= x"C86A0004";
end if;
if first_state_sram_input_id = 8427 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 8428 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 8429 then
	sram_write <= x"C8480008";
end if;
if first_state_sram_input_id = 8430 then
	sram_write <= x"C86A0008";
end if;
if first_state_sram_input_id = 8431 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 8432 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 8433 then
	sram_write <= x"C43C0024";
end if;
if first_state_sram_input_id = 8434 then
	sram_write <= x"8E20841C";
end if;
if first_state_sram_input_id = 8435 then
	sram_write <= x"C8400018";
end if;
if first_state_sram_input_id = 8436 then
	sram_write <= x"C45C0028";
end if;
if first_state_sram_input_id = 8437 then
	sram_write <= x"CC3C0030";
end if;
if first_state_sram_input_id = 8438 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 8439 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 8440 then
	sram_write <= x"03DC0040";
end if;
if first_state_sram_input_id = 8441 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 8442 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 8443 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 8444 then
	sram_write <= x"07DC0040";
end if;
if first_state_sram_input_id = 8445 then
	sram_write <= x"C85C0030";
end if;
if first_state_sram_input_id = 8446 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 8447 then
	sram_write <= x"C03C0028";
end if;
if first_state_sram_input_id = 8448 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 8449 then
	sram_write <= x"03DC0040";
end if;
if first_state_sram_input_id = 8450 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 8451 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 8452 then
	sram_write <= x"82008034";
end if;
if first_state_sram_input_id = 8453 then
	sram_write <= x"07DC0040";
end if;
if first_state_sram_input_id = 8454 then
	sram_write <= x"82008474";
end if;
if first_state_sram_input_id = 8455 then
	sram_write <= x"02420001";
end if;
if first_state_sram_input_id = 8456 then
	sram_write <= x"22440220";
end if;
if first_state_sram_input_id = 8457 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 8458 then
	sram_write <= x"C8400014";
end if;
if first_state_sram_input_id = 8459 then
	sram_write <= x"C45C0038";
end if;
if first_state_sram_input_id = 8460 then
	sram_write <= x"CC3C0030";
end if;
if first_state_sram_input_id = 8461 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 8462 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 8463 then
	sram_write <= x"03DC0044";
end if;
if first_state_sram_input_id = 8464 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 8465 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 8466 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 8467 then
	sram_write <= x"07DC0044";
end if;
if first_state_sram_input_id = 8468 then
	sram_write <= x"C85C0030";
end if;
if first_state_sram_input_id = 8469 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 8470 then
	sram_write <= x"C03C0038";
end if;
if first_state_sram_input_id = 8471 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 8472 then
	sram_write <= x"03DC0044";
end if;
if first_state_sram_input_id = 8473 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 8474 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 8475 then
	sram_write <= x"82008034";
end if;
if first_state_sram_input_id = 8476 then
	sram_write <= x"07DC0044";
end if;
if first_state_sram_input_id = 8477 then
	sram_write <= x"C03C0024";
end if;
if first_state_sram_input_id = 8478 then
	sram_write <= x"06820002";
end if;
if first_state_sram_input_id = 8479 then
	sram_write <= x"C03C0008";
end if;
if first_state_sram_input_id = 8480 then
	sram_write <= x"C05C0004";
end if;
if first_state_sram_input_id = 8481 then
	sram_write <= x"C07C0000";
end if;
if first_state_sram_input_id = 8482 then
	sram_write <= x"82008280";
end if;
if first_state_sram_input_id = 8483 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 8484 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 8485 then
	sram_write <= x"C45C0000";
end if;
if first_state_sram_input_id = 8486 then
	sram_write <= x"C47C0004";
end if;
if first_state_sram_input_id = 8487 then
	sram_write <= x"C43C0008";
end if;
if first_state_sram_input_id = 8488 then
	sram_write <= x"82208524";
end if;
if first_state_sram_input_id = 8489 then
	sram_write <= x"02800354";
end if;
if first_state_sram_input_id = 8490 then
	sram_write <= x"C0880000";
end if;
if first_state_sram_input_id = 8491 then
	sram_write <= x"02A00318";
end if;
if first_state_sram_input_id = 8492 then
	sram_write <= x"C8260000";
end if;
if first_state_sram_input_id = 8493 then
	sram_write <= x"CC2A0000";
end if;
if first_state_sram_input_id = 8494 then
	sram_write <= x"C8260004";
end if;
if first_state_sram_input_id = 8495 then
	sram_write <= x"CC2A0004";
end if;
if first_state_sram_input_id = 8496 then
	sram_write <= x"C8260008";
end if;
if first_state_sram_input_id = 8497 then
	sram_write <= x"CC2A0008";
end if;
if first_state_sram_input_id = 8498 then
	sram_write <= x"02A000C4";
end if;
if first_state_sram_input_id = 8499 then
	sram_write <= x"C0AA0000";
end if;
if first_state_sram_input_id = 8500 then
	sram_write <= x"06AA0001";
end if;
if first_state_sram_input_id = 8501 then
	sram_write <= x"C49C000C";
end if;
if first_state_sram_input_id = 8502 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 8503 then
	sram_write <= x"004A0000";
end if;
if first_state_sram_input_id = 8504 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 8505 then
	sram_write <= x"03DC0018";
end if;
if first_state_sram_input_id = 8506 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 8507 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 8508 then
	sram_write <= x"8200462C";
end if;
if first_state_sram_input_id = 8509 then
	sram_write <= x"07DC0018";
end if;
if first_state_sram_input_id = 8510 then
	sram_write <= x"02800076";
end if;
if first_state_sram_input_id = 8511 then
	sram_write <= x"C03C000C";
end if;
if first_state_sram_input_id = 8512 then
	sram_write <= x"C05C0000";
end if;
if first_state_sram_input_id = 8513 then
	sram_write <= x"C07C0004";
end if;
if first_state_sram_input_id = 8514 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 8515 then
	sram_write <= x"03DC0018";
end if;
if first_state_sram_input_id = 8516 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 8517 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 8518 then
	sram_write <= x"82008280";
end if;
if first_state_sram_input_id = 8519 then
	sram_write <= x"07DC0018";
end if;
if first_state_sram_input_id = 8520 then
	sram_write <= x"82008524";
end if;
if first_state_sram_input_id = 8521 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 8522 then
	sram_write <= x"C05C0008";
end if;
if first_state_sram_input_id = 8523 then
	sram_write <= x"824285B4";
end if;
if first_state_sram_input_id = 8524 then
	sram_write <= x"02200354";
end if;
if first_state_sram_input_id = 8525 then
	sram_write <= x"C0220004";
end if;
if first_state_sram_input_id = 8526 then
	sram_write <= x"02600318";
end if;
if first_state_sram_input_id = 8527 then
	sram_write <= x"C09C0004";
end if;
if first_state_sram_input_id = 8528 then
	sram_write <= x"C8280000";
end if;
if first_state_sram_input_id = 8529 then
	sram_write <= x"CC260000";
end if;
if first_state_sram_input_id = 8530 then
	sram_write <= x"C8280004";
end if;
if first_state_sram_input_id = 8531 then
	sram_write <= x"CC260004";
end if;
if first_state_sram_input_id = 8532 then
	sram_write <= x"C8280008";
end if;
if first_state_sram_input_id = 8533 then
	sram_write <= x"CC260008";
end if;
if first_state_sram_input_id = 8534 then
	sram_write <= x"026000C4";
end if;
if first_state_sram_input_id = 8535 then
	sram_write <= x"C0660000";
end if;
if first_state_sram_input_id = 8536 then
	sram_write <= x"06660001";
end if;
if first_state_sram_input_id = 8537 then
	sram_write <= x"C43C0010";
end if;
if first_state_sram_input_id = 8538 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 8539 then
	sram_write <= x"00460000";
end if;
if first_state_sram_input_id = 8540 then
	sram_write <= x"00280000";
end if;
if first_state_sram_input_id = 8541 then
	sram_write <= x"03DC001C";
end if;
if first_state_sram_input_id = 8542 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 8543 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 8544 then
	sram_write <= x"8200462C";
end if;
if first_state_sram_input_id = 8545 then
	sram_write <= x"07DC001C";
end if;
if first_state_sram_input_id = 8546 then
	sram_write <= x"02800076";
end if;
if first_state_sram_input_id = 8547 then
	sram_write <= x"C03C0010";
end if;
if first_state_sram_input_id = 8548 then
	sram_write <= x"C05C0000";
end if;
if first_state_sram_input_id = 8549 then
	sram_write <= x"C07C0004";
end if;
if first_state_sram_input_id = 8550 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 8551 then
	sram_write <= x"03DC001C";
end if;
if first_state_sram_input_id = 8552 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 8553 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 8554 then
	sram_write <= x"82008280";
end if;
if first_state_sram_input_id = 8555 then
	sram_write <= x"07DC001C";
end if;
if first_state_sram_input_id = 8556 then
	sram_write <= x"820085B4";
end if;
if first_state_sram_input_id = 8557 then
	sram_write <= x"02200002";
end if;
if first_state_sram_input_id = 8558 then
	sram_write <= x"C05C0008";
end if;
if first_state_sram_input_id = 8559 then
	sram_write <= x"82428644";
end if;
if first_state_sram_input_id = 8560 then
	sram_write <= x"02200354";
end if;
if first_state_sram_input_id = 8561 then
	sram_write <= x"C0220008";
end if;
if first_state_sram_input_id = 8562 then
	sram_write <= x"02600318";
end if;
if first_state_sram_input_id = 8563 then
	sram_write <= x"C09C0004";
end if;
if first_state_sram_input_id = 8564 then
	sram_write <= x"C8280000";
end if;
if first_state_sram_input_id = 8565 then
	sram_write <= x"CC260000";
end if;
if first_state_sram_input_id = 8566 then
	sram_write <= x"C8280004";
end if;
if first_state_sram_input_id = 8567 then
	sram_write <= x"CC260004";
end if;
if first_state_sram_input_id = 8568 then
	sram_write <= x"C8280008";
end if;
if first_state_sram_input_id = 8569 then
	sram_write <= x"CC260008";
end if;
if first_state_sram_input_id = 8570 then
	sram_write <= x"026000C4";
end if;
if first_state_sram_input_id = 8571 then
	sram_write <= x"C0660000";
end if;
if first_state_sram_input_id = 8572 then
	sram_write <= x"06660001";
end if;
if first_state_sram_input_id = 8573 then
	sram_write <= x"C43C0014";
end if;
if first_state_sram_input_id = 8574 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 8575 then
	sram_write <= x"00460000";
end if;
if first_state_sram_input_id = 8576 then
	sram_write <= x"00280000";
end if;
if first_state_sram_input_id = 8577 then
	sram_write <= x"03DC0020";
end if;
if first_state_sram_input_id = 8578 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 8579 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 8580 then
	sram_write <= x"8200462C";
end if;
if first_state_sram_input_id = 8581 then
	sram_write <= x"07DC0020";
end if;
if first_state_sram_input_id = 8582 then
	sram_write <= x"02800076";
end if;
if first_state_sram_input_id = 8583 then
	sram_write <= x"C03C0014";
end if;
if first_state_sram_input_id = 8584 then
	sram_write <= x"C05C0000";
end if;
if first_state_sram_input_id = 8585 then
	sram_write <= x"C07C0004";
end if;
if first_state_sram_input_id = 8586 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 8587 then
	sram_write <= x"03DC0020";
end if;
if first_state_sram_input_id = 8588 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 8589 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 8590 then
	sram_write <= x"82008280";
end if;
if first_state_sram_input_id = 8591 then
	sram_write <= x"07DC0020";
end if;
if first_state_sram_input_id = 8592 then
	sram_write <= x"82008644";
end if;
if first_state_sram_input_id = 8593 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 8594 then
	sram_write <= x"C05C0008";
end if;
if first_state_sram_input_id = 8595 then
	sram_write <= x"824286D4";
end if;
if first_state_sram_input_id = 8596 then
	sram_write <= x"02200354";
end if;
if first_state_sram_input_id = 8597 then
	sram_write <= x"C022000C";
end if;
if first_state_sram_input_id = 8598 then
	sram_write <= x"02600318";
end if;
if first_state_sram_input_id = 8599 then
	sram_write <= x"C09C0004";
end if;
if first_state_sram_input_id = 8600 then
	sram_write <= x"C8280000";
end if;
if first_state_sram_input_id = 8601 then
	sram_write <= x"CC260000";
end if;
if first_state_sram_input_id = 8602 then
	sram_write <= x"C8280004";
end if;
if first_state_sram_input_id = 8603 then
	sram_write <= x"CC260004";
end if;
if first_state_sram_input_id = 8604 then
	sram_write <= x"C8280008";
end if;
if first_state_sram_input_id = 8605 then
	sram_write <= x"CC260008";
end if;
if first_state_sram_input_id = 8606 then
	sram_write <= x"026000C4";
end if;
if first_state_sram_input_id = 8607 then
	sram_write <= x"C0660000";
end if;
if first_state_sram_input_id = 8608 then
	sram_write <= x"06660001";
end if;
if first_state_sram_input_id = 8609 then
	sram_write <= x"C43C0018";
end if;
if first_state_sram_input_id = 8610 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 8611 then
	sram_write <= x"00460000";
end if;
if first_state_sram_input_id = 8612 then
	sram_write <= x"00280000";
end if;
if first_state_sram_input_id = 8613 then
	sram_write <= x"03DC0024";
end if;
if first_state_sram_input_id = 8614 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 8615 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 8616 then
	sram_write <= x"8200462C";
end if;
if first_state_sram_input_id = 8617 then
	sram_write <= x"07DC0024";
end if;
if first_state_sram_input_id = 8618 then
	sram_write <= x"02800076";
end if;
if first_state_sram_input_id = 8619 then
	sram_write <= x"C03C0018";
end if;
if first_state_sram_input_id = 8620 then
	sram_write <= x"C05C0000";
end if;
if first_state_sram_input_id = 8621 then
	sram_write <= x"C07C0004";
end if;
if first_state_sram_input_id = 8622 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 8623 then
	sram_write <= x"03DC0024";
end if;
if first_state_sram_input_id = 8624 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 8625 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 8626 then
	sram_write <= x"82008280";
end if;
if first_state_sram_input_id = 8627 then
	sram_write <= x"07DC0024";
end if;
if first_state_sram_input_id = 8628 then
	sram_write <= x"820086D4";
end if;
if first_state_sram_input_id = 8629 then
	sram_write <= x"02200004";
end if;
if first_state_sram_input_id = 8630 then
	sram_write <= x"C05C0008";
end if;
if first_state_sram_input_id = 8631 then
	sram_write <= x"82428748";
end if;
if first_state_sram_input_id = 8632 then
	sram_write <= x"02200354";
end if;
if first_state_sram_input_id = 8633 then
	sram_write <= x"C0220010";
end if;
if first_state_sram_input_id = 8634 then
	sram_write <= x"02400318";
end if;
if first_state_sram_input_id = 8635 then
	sram_write <= x"C07C0004";
end if;
if first_state_sram_input_id = 8636 then
	sram_write <= x"C8260000";
end if;
if first_state_sram_input_id = 8637 then
	sram_write <= x"CC240000";
end if;
if first_state_sram_input_id = 8638 then
	sram_write <= x"C8260004";
end if;
if first_state_sram_input_id = 8639 then
	sram_write <= x"CC240004";
end if;
if first_state_sram_input_id = 8640 then
	sram_write <= x"C8260008";
end if;
if first_state_sram_input_id = 8641 then
	sram_write <= x"CC240008";
end if;
if first_state_sram_input_id = 8642 then
	sram_write <= x"024000C4";
end if;
if first_state_sram_input_id = 8643 then
	sram_write <= x"C0440000";
end if;
if first_state_sram_input_id = 8644 then
	sram_write <= x"06440001";
end if;
if first_state_sram_input_id = 8645 then
	sram_write <= x"C43C001C";
end if;
if first_state_sram_input_id = 8646 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 8647 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 8648 then
	sram_write <= x"03DC0028";
end if;
if first_state_sram_input_id = 8649 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 8650 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 8651 then
	sram_write <= x"8200462C";
end if;
if first_state_sram_input_id = 8652 then
	sram_write <= x"07DC0028";
end if;
if first_state_sram_input_id = 8653 then
	sram_write <= x"02800076";
end if;
if first_state_sram_input_id = 8654 then
	sram_write <= x"C03C001C";
end if;
if first_state_sram_input_id = 8655 then
	sram_write <= x"C05C0000";
end if;
if first_state_sram_input_id = 8656 then
	sram_write <= x"C07C0004";
end if;
if first_state_sram_input_id = 8657 then
	sram_write <= x"82008280";
end if;
if first_state_sram_input_id = 8658 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 8659 then
	sram_write <= x"C0620014";
end if;
if first_state_sram_input_id = 8660 then
	sram_write <= x"C082001C";
end if;
if first_state_sram_input_id = 8661 then
	sram_write <= x"C0A20004";
end if;
if first_state_sram_input_id = 8662 then
	sram_write <= x"C0C20010";
end if;
if first_state_sram_input_id = 8663 then
	sram_write <= x"02E002E0";
end if;
if first_state_sram_input_id = 8664 then
	sram_write <= x"23040220";
end if;
if first_state_sram_input_id = 8665 then
	sram_write <= x"D0670000";
end if;
if first_state_sram_input_id = 8666 then
	sram_write <= x"C8260000";
end if;
if first_state_sram_input_id = 8667 then
	sram_write <= x"CC2E0000";
end if;
if first_state_sram_input_id = 8668 then
	sram_write <= x"C8260004";
end if;
if first_state_sram_input_id = 8669 then
	sram_write <= x"CC2E0004";
end if;
if first_state_sram_input_id = 8670 then
	sram_write <= x"C8260008";
end if;
if first_state_sram_input_id = 8671 then
	sram_write <= x"CC2E0008";
end if;
if first_state_sram_input_id = 8672 then
	sram_write <= x"C0220018";
end if;
if first_state_sram_input_id = 8673 then
	sram_write <= x"C0220000";
end if;
if first_state_sram_input_id = 8674 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 8675 then
	sram_write <= x"D0686000";
end if;
if first_state_sram_input_id = 8676 then
	sram_write <= x"22840220";
end if;
if first_state_sram_input_id = 8677 then
	sram_write <= x"D08A8000";
end if;
if first_state_sram_input_id = 8678 then
	sram_write <= x"C4FC0000";
end if;
if first_state_sram_input_id = 8679 then
	sram_write <= x"C4DC0004";
end if;
if first_state_sram_input_id = 8680 then
	sram_write <= x"C45C0008";
end if;
if first_state_sram_input_id = 8681 then
	sram_write <= x"C47C000C";
end if;
if first_state_sram_input_id = 8682 then
	sram_write <= x"C49C0010";
end if;
if first_state_sram_input_id = 8683 then
	sram_write <= x"C43C0014";
end if;
if first_state_sram_input_id = 8684 then
	sram_write <= x"82208914";
end if;
if first_state_sram_input_id = 8685 then
	sram_write <= x"02A00354";
end if;
if first_state_sram_input_id = 8686 then
	sram_write <= x"C0AA0000";
end if;
if first_state_sram_input_id = 8687 then
	sram_write <= x"03000318";
end if;
if first_state_sram_input_id = 8688 then
	sram_write <= x"C8280000";
end if;
if first_state_sram_input_id = 8689 then
	sram_write <= x"CC300000";
end if;
if first_state_sram_input_id = 8690 then
	sram_write <= x"C8280004";
end if;
if first_state_sram_input_id = 8691 then
	sram_write <= x"CC300004";
end if;
if first_state_sram_input_id = 8692 then
	sram_write <= x"C8280008";
end if;
if first_state_sram_input_id = 8693 then
	sram_write <= x"CC300008";
end if;
if first_state_sram_input_id = 8694 then
	sram_write <= x"030000C4";
end if;
if first_state_sram_input_id = 8695 then
	sram_write <= x"C1100000";
end if;
if first_state_sram_input_id = 8696 then
	sram_write <= x"07100001";
end if;
if first_state_sram_input_id = 8697 then
	sram_write <= x"C4BC0018";
end if;
if first_state_sram_input_id = 8698 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 8699 then
	sram_write <= x"00500000";
end if;
if first_state_sram_input_id = 8700 then
	sram_write <= x"00280000";
end if;
if first_state_sram_input_id = 8701 then
	sram_write <= x"03DC0024";
end if;
if first_state_sram_input_id = 8702 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 8703 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 8704 then
	sram_write <= x"8200462C";
end if;
if first_state_sram_input_id = 8705 then
	sram_write <= x"07DC0024";
end if;
if first_state_sram_input_id = 8706 then
	sram_write <= x"C03C0018";
end if;
if first_state_sram_input_id = 8707 then
	sram_write <= x"C04201D8";
end if;
if first_state_sram_input_id = 8708 then
	sram_write <= x"C0640000";
end if;
if first_state_sram_input_id = 8709 then
	sram_write <= x"C8260000";
end if;
if first_state_sram_input_id = 8710 then
	sram_write <= x"C09C000C";
end if;
if first_state_sram_input_id = 8711 then
	sram_write <= x"C8480000";
end if;
if first_state_sram_input_id = 8712 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 8713 then
	sram_write <= x"C8460004";
end if;
if first_state_sram_input_id = 8714 then
	sram_write <= x"C8680004";
end if;
if first_state_sram_input_id = 8715 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 8716 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 8717 then
	sram_write <= x"C8460008";
end if;
if first_state_sram_input_id = 8718 then
	sram_write <= x"C8680008";
end if;
if first_state_sram_input_id = 8719 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 8720 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 8721 then
	sram_write <= x"8E208898";
end if;
if first_state_sram_input_id = 8722 then
	sram_write <= x"C8400018";
end if;
if first_state_sram_input_id = 8723 then
	sram_write <= x"C45C001C";
end if;
if first_state_sram_input_id = 8724 then
	sram_write <= x"CC3C0020";
end if;
if first_state_sram_input_id = 8725 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 8726 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 8727 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 8728 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 8729 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 8730 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 8731 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 8732 then
	sram_write <= x"C85C0020";
end if;
if first_state_sram_input_id = 8733 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 8734 then
	sram_write <= x"C03C001C";
end if;
if first_state_sram_input_id = 8735 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 8736 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 8737 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 8738 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 8739 then
	sram_write <= x"82008034";
end if;
if first_state_sram_input_id = 8740 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 8741 then
	sram_write <= x"820088E8";
end if;
if first_state_sram_input_id = 8742 then
	sram_write <= x"C04201DC";
end if;
if first_state_sram_input_id = 8743 then
	sram_write <= x"C8400014";
end if;
if first_state_sram_input_id = 8744 then
	sram_write <= x"C45C0028";
end if;
if first_state_sram_input_id = 8745 then
	sram_write <= x"CC3C0020";
end if;
if first_state_sram_input_id = 8746 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 8747 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 8748 then
	sram_write <= x"03DC0034";
end if;
if first_state_sram_input_id = 8749 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 8750 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 8751 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 8752 then
	sram_write <= x"07DC0034";
end if;
if first_state_sram_input_id = 8753 then
	sram_write <= x"C85C0020";
end if;
if first_state_sram_input_id = 8754 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 8755 then
	sram_write <= x"C03C0028";
end if;
if first_state_sram_input_id = 8756 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 8757 then
	sram_write <= x"03DC0034";
end if;
if first_state_sram_input_id = 8758 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 8759 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 8760 then
	sram_write <= x"82008034";
end if;
if first_state_sram_input_id = 8761 then
	sram_write <= x"07DC0034";
end if;
if first_state_sram_input_id = 8762 then
	sram_write <= x"02800074";
end if;
if first_state_sram_input_id = 8763 then
	sram_write <= x"C03C0018";
end if;
if first_state_sram_input_id = 8764 then
	sram_write <= x"C05C000C";
end if;
if first_state_sram_input_id = 8765 then
	sram_write <= x"C07C0010";
end if;
if first_state_sram_input_id = 8766 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 8767 then
	sram_write <= x"03DC0034";
end if;
if first_state_sram_input_id = 8768 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 8769 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 8770 then
	sram_write <= x"82008280";
end if;
if first_state_sram_input_id = 8771 then
	sram_write <= x"07DC0034";
end if;
if first_state_sram_input_id = 8772 then
	sram_write <= x"82008914";
end if;
if first_state_sram_input_id = 8773 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 8774 then
	sram_write <= x"C05C0014";
end if;
if first_state_sram_input_id = 8775 then
	sram_write <= x"82428A84";
end if;
if first_state_sram_input_id = 8776 then
	sram_write <= x"02200354";
end if;
if first_state_sram_input_id = 8777 then
	sram_write <= x"C0220004";
end if;
if first_state_sram_input_id = 8778 then
	sram_write <= x"02600318";
end if;
if first_state_sram_input_id = 8779 then
	sram_write <= x"C09C0010";
end if;
if first_state_sram_input_id = 8780 then
	sram_write <= x"C8280000";
end if;
if first_state_sram_input_id = 8781 then
	sram_write <= x"CC260000";
end if;
if first_state_sram_input_id = 8782 then
	sram_write <= x"C8280004";
end if;
if first_state_sram_input_id = 8783 then
	sram_write <= x"CC260004";
end if;
if first_state_sram_input_id = 8784 then
	sram_write <= x"C8280008";
end if;
if first_state_sram_input_id = 8785 then
	sram_write <= x"CC260008";
end if;
if first_state_sram_input_id = 8786 then
	sram_write <= x"026000C4";
end if;
if first_state_sram_input_id = 8787 then
	sram_write <= x"C0660000";
end if;
if first_state_sram_input_id = 8788 then
	sram_write <= x"06660001";
end if;
if first_state_sram_input_id = 8789 then
	sram_write <= x"C43C002C";
end if;
if first_state_sram_input_id = 8790 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 8791 then
	sram_write <= x"00460000";
end if;
if first_state_sram_input_id = 8792 then
	sram_write <= x"00280000";
end if;
if first_state_sram_input_id = 8793 then
	sram_write <= x"03DC0038";
end if;
if first_state_sram_input_id = 8794 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 8795 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 8796 then
	sram_write <= x"8200462C";
end if;
if first_state_sram_input_id = 8797 then
	sram_write <= x"07DC0038";
end if;
if first_state_sram_input_id = 8798 then
	sram_write <= x"C03C002C";
end if;
if first_state_sram_input_id = 8799 then
	sram_write <= x"C04201D8";
end if;
if first_state_sram_input_id = 8800 then
	sram_write <= x"C0640000";
end if;
if first_state_sram_input_id = 8801 then
	sram_write <= x"C8260000";
end if;
if first_state_sram_input_id = 8802 then
	sram_write <= x"C09C000C";
end if;
if first_state_sram_input_id = 8803 then
	sram_write <= x"C8480000";
end if;
if first_state_sram_input_id = 8804 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 8805 then
	sram_write <= x"C8460004";
end if;
if first_state_sram_input_id = 8806 then
	sram_write <= x"C8680004";
end if;
if first_state_sram_input_id = 8807 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 8808 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 8809 then
	sram_write <= x"C8460008";
end if;
if first_state_sram_input_id = 8810 then
	sram_write <= x"C8680008";
end if;
if first_state_sram_input_id = 8811 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 8812 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 8813 then
	sram_write <= x"8E208A08";
end if;
if first_state_sram_input_id = 8814 then
	sram_write <= x"C8400018";
end if;
if first_state_sram_input_id = 8815 then
	sram_write <= x"C45C0030";
end if;
if first_state_sram_input_id = 8816 then
	sram_write <= x"CC3C0038";
end if;
if first_state_sram_input_id = 8817 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 8818 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 8819 then
	sram_write <= x"03DC0048";
end if;
if first_state_sram_input_id = 8820 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 8821 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 8822 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 8823 then
	sram_write <= x"07DC0048";
end if;
if first_state_sram_input_id = 8824 then
	sram_write <= x"C85C0038";
end if;
if first_state_sram_input_id = 8825 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 8826 then
	sram_write <= x"C03C0030";
end if;
if first_state_sram_input_id = 8827 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 8828 then
	sram_write <= x"03DC0048";
end if;
if first_state_sram_input_id = 8829 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 8830 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 8831 then
	sram_write <= x"82008034";
end if;
if first_state_sram_input_id = 8832 then
	sram_write <= x"07DC0048";
end if;
if first_state_sram_input_id = 8833 then
	sram_write <= x"82008A58";
end if;
if first_state_sram_input_id = 8834 then
	sram_write <= x"C04201DC";
end if;
if first_state_sram_input_id = 8835 then
	sram_write <= x"C8400014";
end if;
if first_state_sram_input_id = 8836 then
	sram_write <= x"C45C0040";
end if;
if first_state_sram_input_id = 8837 then
	sram_write <= x"CC3C0038";
end if;
if first_state_sram_input_id = 8838 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 8839 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 8840 then
	sram_write <= x"03DC004C";
end if;
if first_state_sram_input_id = 8841 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 8842 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 8843 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 8844 then
	sram_write <= x"07DC004C";
end if;
if first_state_sram_input_id = 8845 then
	sram_write <= x"C85C0038";
end if;
if first_state_sram_input_id = 8846 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 8847 then
	sram_write <= x"C03C0040";
end if;
if first_state_sram_input_id = 8848 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 8849 then
	sram_write <= x"03DC004C";
end if;
if first_state_sram_input_id = 8850 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 8851 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 8852 then
	sram_write <= x"82008034";
end if;
if first_state_sram_input_id = 8853 then
	sram_write <= x"07DC004C";
end if;
if first_state_sram_input_id = 8854 then
	sram_write <= x"02800074";
end if;
if first_state_sram_input_id = 8855 then
	sram_write <= x"C03C002C";
end if;
if first_state_sram_input_id = 8856 then
	sram_write <= x"C05C000C";
end if;
if first_state_sram_input_id = 8857 then
	sram_write <= x"C07C0010";
end if;
if first_state_sram_input_id = 8858 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 8859 then
	sram_write <= x"03DC004C";
end if;
if first_state_sram_input_id = 8860 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 8861 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 8862 then
	sram_write <= x"82008280";
end if;
if first_state_sram_input_id = 8863 then
	sram_write <= x"07DC004C";
end if;
if first_state_sram_input_id = 8864 then
	sram_write <= x"82008A84";
end if;
if first_state_sram_input_id = 8865 then
	sram_write <= x"02200002";
end if;
if first_state_sram_input_id = 8866 then
	sram_write <= x"C05C0014";
end if;
if first_state_sram_input_id = 8867 then
	sram_write <= x"82428BF4";
end if;
if first_state_sram_input_id = 8868 then
	sram_write <= x"02200354";
end if;
if first_state_sram_input_id = 8869 then
	sram_write <= x"C0220008";
end if;
if first_state_sram_input_id = 8870 then
	sram_write <= x"02600318";
end if;
if first_state_sram_input_id = 8871 then
	sram_write <= x"C09C0010";
end if;
if first_state_sram_input_id = 8872 then
	sram_write <= x"C8280000";
end if;
if first_state_sram_input_id = 8873 then
	sram_write <= x"CC260000";
end if;
if first_state_sram_input_id = 8874 then
	sram_write <= x"C8280004";
end if;
if first_state_sram_input_id = 8875 then
	sram_write <= x"CC260004";
end if;
if first_state_sram_input_id = 8876 then
	sram_write <= x"C8280008";
end if;
if first_state_sram_input_id = 8877 then
	sram_write <= x"CC260008";
end if;
if first_state_sram_input_id = 8878 then
	sram_write <= x"026000C4";
end if;
if first_state_sram_input_id = 8879 then
	sram_write <= x"C0660000";
end if;
if first_state_sram_input_id = 8880 then
	sram_write <= x"06660001";
end if;
if first_state_sram_input_id = 8881 then
	sram_write <= x"C43C0044";
end if;
if first_state_sram_input_id = 8882 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 8883 then
	sram_write <= x"00460000";
end if;
if first_state_sram_input_id = 8884 then
	sram_write <= x"00280000";
end if;
if first_state_sram_input_id = 8885 then
	sram_write <= x"03DC0050";
end if;
if first_state_sram_input_id = 8886 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 8887 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 8888 then
	sram_write <= x"8200462C";
end if;
if first_state_sram_input_id = 8889 then
	sram_write <= x"07DC0050";
end if;
if first_state_sram_input_id = 8890 then
	sram_write <= x"C03C0044";
end if;
if first_state_sram_input_id = 8891 then
	sram_write <= x"C04201D8";
end if;
if first_state_sram_input_id = 8892 then
	sram_write <= x"C0640000";
end if;
if first_state_sram_input_id = 8893 then
	sram_write <= x"C8260000";
end if;
if first_state_sram_input_id = 8894 then
	sram_write <= x"C09C000C";
end if;
if first_state_sram_input_id = 8895 then
	sram_write <= x"C8480000";
end if;
if first_state_sram_input_id = 8896 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 8897 then
	sram_write <= x"C8460004";
end if;
if first_state_sram_input_id = 8898 then
	sram_write <= x"C8680004";
end if;
if first_state_sram_input_id = 8899 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 8900 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 8901 then
	sram_write <= x"C8460008";
end if;
if first_state_sram_input_id = 8902 then
	sram_write <= x"C8680008";
end if;
if first_state_sram_input_id = 8903 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 8904 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 8905 then
	sram_write <= x"8E208B78";
end if;
if first_state_sram_input_id = 8906 then
	sram_write <= x"C8400018";
end if;
if first_state_sram_input_id = 8907 then
	sram_write <= x"C45C0048";
end if;
if first_state_sram_input_id = 8908 then
	sram_write <= x"CC3C0050";
end if;
if first_state_sram_input_id = 8909 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 8910 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 8911 then
	sram_write <= x"03DC0060";
end if;
if first_state_sram_input_id = 8912 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 8913 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 8914 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 8915 then
	sram_write <= x"07DC0060";
end if;
if first_state_sram_input_id = 8916 then
	sram_write <= x"C85C0050";
end if;
if first_state_sram_input_id = 8917 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 8918 then
	sram_write <= x"C03C0048";
end if;
if first_state_sram_input_id = 8919 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 8920 then
	sram_write <= x"03DC0060";
end if;
if first_state_sram_input_id = 8921 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 8922 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 8923 then
	sram_write <= x"82008034";
end if;
if first_state_sram_input_id = 8924 then
	sram_write <= x"07DC0060";
end if;
if first_state_sram_input_id = 8925 then
	sram_write <= x"82008BC8";
end if;
if first_state_sram_input_id = 8926 then
	sram_write <= x"C04201DC";
end if;
if first_state_sram_input_id = 8927 then
	sram_write <= x"C8400014";
end if;
if first_state_sram_input_id = 8928 then
	sram_write <= x"C45C0058";
end if;
if first_state_sram_input_id = 8929 then
	sram_write <= x"CC3C0050";
end if;
if first_state_sram_input_id = 8930 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 8931 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 8932 then
	sram_write <= x"03DC0064";
end if;
if first_state_sram_input_id = 8933 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 8934 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 8935 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 8936 then
	sram_write <= x"07DC0064";
end if;
if first_state_sram_input_id = 8937 then
	sram_write <= x"C85C0050";
end if;
if first_state_sram_input_id = 8938 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 8939 then
	sram_write <= x"C03C0058";
end if;
if first_state_sram_input_id = 8940 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 8941 then
	sram_write <= x"03DC0064";
end if;
if first_state_sram_input_id = 8942 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 8943 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 8944 then
	sram_write <= x"82008034";
end if;
if first_state_sram_input_id = 8945 then
	sram_write <= x"07DC0064";
end if;
if first_state_sram_input_id = 8946 then
	sram_write <= x"02800074";
end if;
if first_state_sram_input_id = 8947 then
	sram_write <= x"C03C0044";
end if;
if first_state_sram_input_id = 8948 then
	sram_write <= x"C05C000C";
end if;
if first_state_sram_input_id = 8949 then
	sram_write <= x"C07C0010";
end if;
if first_state_sram_input_id = 8950 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 8951 then
	sram_write <= x"03DC0064";
end if;
if first_state_sram_input_id = 8952 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 8953 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 8954 then
	sram_write <= x"82008280";
end if;
if first_state_sram_input_id = 8955 then
	sram_write <= x"07DC0064";
end if;
if first_state_sram_input_id = 8956 then
	sram_write <= x"82008BF4";
end if;
if first_state_sram_input_id = 8957 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 8958 then
	sram_write <= x"C05C0014";
end if;
if first_state_sram_input_id = 8959 then
	sram_write <= x"82428D64";
end if;
if first_state_sram_input_id = 8960 then
	sram_write <= x"02200354";
end if;
if first_state_sram_input_id = 8961 then
	sram_write <= x"C022000C";
end if;
if first_state_sram_input_id = 8962 then
	sram_write <= x"02600318";
end if;
if first_state_sram_input_id = 8963 then
	sram_write <= x"C09C0010";
end if;
if first_state_sram_input_id = 8964 then
	sram_write <= x"C8280000";
end if;
if first_state_sram_input_id = 8965 then
	sram_write <= x"CC260000";
end if;
if first_state_sram_input_id = 8966 then
	sram_write <= x"C8280004";
end if;
if first_state_sram_input_id = 8967 then
	sram_write <= x"CC260004";
end if;
if first_state_sram_input_id = 8968 then
	sram_write <= x"C8280008";
end if;
if first_state_sram_input_id = 8969 then
	sram_write <= x"CC260008";
end if;
if first_state_sram_input_id = 8970 then
	sram_write <= x"026000C4";
end if;
if first_state_sram_input_id = 8971 then
	sram_write <= x"C0660000";
end if;
if first_state_sram_input_id = 8972 then
	sram_write <= x"06660001";
end if;
if first_state_sram_input_id = 8973 then
	sram_write <= x"C43C005C";
end if;
if first_state_sram_input_id = 8974 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 8975 then
	sram_write <= x"00460000";
end if;
if first_state_sram_input_id = 8976 then
	sram_write <= x"00280000";
end if;
if first_state_sram_input_id = 8977 then
	sram_write <= x"03DC0068";
end if;
if first_state_sram_input_id = 8978 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 8979 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 8980 then
	sram_write <= x"8200462C";
end if;
if first_state_sram_input_id = 8981 then
	sram_write <= x"07DC0068";
end if;
if first_state_sram_input_id = 8982 then
	sram_write <= x"C03C005C";
end if;
if first_state_sram_input_id = 8983 then
	sram_write <= x"C04201D8";
end if;
if first_state_sram_input_id = 8984 then
	sram_write <= x"C0640000";
end if;
if first_state_sram_input_id = 8985 then
	sram_write <= x"C8260000";
end if;
if first_state_sram_input_id = 8986 then
	sram_write <= x"C09C000C";
end if;
if first_state_sram_input_id = 8987 then
	sram_write <= x"C8480000";
end if;
if first_state_sram_input_id = 8988 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 8989 then
	sram_write <= x"C8460004";
end if;
if first_state_sram_input_id = 8990 then
	sram_write <= x"C8680004";
end if;
if first_state_sram_input_id = 8991 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 8992 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 8993 then
	sram_write <= x"C8460008";
end if;
if first_state_sram_input_id = 8994 then
	sram_write <= x"C8680008";
end if;
if first_state_sram_input_id = 8995 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 8996 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 8997 then
	sram_write <= x"8E208CE8";
end if;
if first_state_sram_input_id = 8998 then
	sram_write <= x"C8400018";
end if;
if first_state_sram_input_id = 8999 then
	sram_write <= x"C45C0060";
end if;
if first_state_sram_input_id = 9000 then
	sram_write <= x"CC3C0068";
end if;
if first_state_sram_input_id = 9001 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 9002 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 9003 then
	sram_write <= x"03DC0078";
end if;
if first_state_sram_input_id = 9004 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 9005 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 9006 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 9007 then
	sram_write <= x"07DC0078";
end if;
if first_state_sram_input_id = 9008 then
	sram_write <= x"C85C0068";
end if;
if first_state_sram_input_id = 9009 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 9010 then
	sram_write <= x"C03C0060";
end if;
if first_state_sram_input_id = 9011 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 9012 then
	sram_write <= x"03DC0078";
end if;
if first_state_sram_input_id = 9013 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 9014 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 9015 then
	sram_write <= x"82008034";
end if;
if first_state_sram_input_id = 9016 then
	sram_write <= x"07DC0078";
end if;
if first_state_sram_input_id = 9017 then
	sram_write <= x"82008D38";
end if;
if first_state_sram_input_id = 9018 then
	sram_write <= x"C04201DC";
end if;
if first_state_sram_input_id = 9019 then
	sram_write <= x"C8400014";
end if;
if first_state_sram_input_id = 9020 then
	sram_write <= x"C45C0070";
end if;
if first_state_sram_input_id = 9021 then
	sram_write <= x"CC3C0068";
end if;
if first_state_sram_input_id = 9022 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 9023 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 9024 then
	sram_write <= x"03DC007C";
end if;
if first_state_sram_input_id = 9025 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 9026 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 9027 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 9028 then
	sram_write <= x"07DC007C";
end if;
if first_state_sram_input_id = 9029 then
	sram_write <= x"C85C0068";
end if;
if first_state_sram_input_id = 9030 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 9031 then
	sram_write <= x"C03C0070";
end if;
if first_state_sram_input_id = 9032 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 9033 then
	sram_write <= x"03DC007C";
end if;
if first_state_sram_input_id = 9034 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 9035 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 9036 then
	sram_write <= x"82008034";
end if;
if first_state_sram_input_id = 9037 then
	sram_write <= x"07DC007C";
end if;
if first_state_sram_input_id = 9038 then
	sram_write <= x"02800074";
end if;
if first_state_sram_input_id = 9039 then
	sram_write <= x"C03C005C";
end if;
if first_state_sram_input_id = 9040 then
	sram_write <= x"C05C000C";
end if;
if first_state_sram_input_id = 9041 then
	sram_write <= x"C07C0010";
end if;
if first_state_sram_input_id = 9042 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 9043 then
	sram_write <= x"03DC007C";
end if;
if first_state_sram_input_id = 9044 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 9045 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 9046 then
	sram_write <= x"82008280";
end if;
if first_state_sram_input_id = 9047 then
	sram_write <= x"07DC007C";
end if;
if first_state_sram_input_id = 9048 then
	sram_write <= x"82008D64";
end if;
if first_state_sram_input_id = 9049 then
	sram_write <= x"02200004";
end if;
if first_state_sram_input_id = 9050 then
	sram_write <= x"C05C0014";
end if;
if first_state_sram_input_id = 9051 then
	sram_write <= x"82428ED0";
end if;
if first_state_sram_input_id = 9052 then
	sram_write <= x"02200354";
end if;
if first_state_sram_input_id = 9053 then
	sram_write <= x"C0220010";
end if;
if first_state_sram_input_id = 9054 then
	sram_write <= x"02400318";
end if;
if first_state_sram_input_id = 9055 then
	sram_write <= x"C07C0010";
end if;
if first_state_sram_input_id = 9056 then
	sram_write <= x"C8260000";
end if;
if first_state_sram_input_id = 9057 then
	sram_write <= x"CC240000";
end if;
if first_state_sram_input_id = 9058 then
	sram_write <= x"C8260004";
end if;
if first_state_sram_input_id = 9059 then
	sram_write <= x"CC240004";
end if;
if first_state_sram_input_id = 9060 then
	sram_write <= x"C8260008";
end if;
if first_state_sram_input_id = 9061 then
	sram_write <= x"CC240008";
end if;
if first_state_sram_input_id = 9062 then
	sram_write <= x"024000C4";
end if;
if first_state_sram_input_id = 9063 then
	sram_write <= x"C0440000";
end if;
if first_state_sram_input_id = 9064 then
	sram_write <= x"06440001";
end if;
if first_state_sram_input_id = 9065 then
	sram_write <= x"C43C0074";
end if;
if first_state_sram_input_id = 9066 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 9067 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 9068 then
	sram_write <= x"03DC0080";
end if;
if first_state_sram_input_id = 9069 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 9070 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 9071 then
	sram_write <= x"8200462C";
end if;
if first_state_sram_input_id = 9072 then
	sram_write <= x"07DC0080";
end if;
if first_state_sram_input_id = 9073 then
	sram_write <= x"C03C0074";
end if;
if first_state_sram_input_id = 9074 then
	sram_write <= x"C04201D8";
end if;
if first_state_sram_input_id = 9075 then
	sram_write <= x"C0640000";
end if;
if first_state_sram_input_id = 9076 then
	sram_write <= x"C8260000";
end if;
if first_state_sram_input_id = 9077 then
	sram_write <= x"C09C000C";
end if;
if first_state_sram_input_id = 9078 then
	sram_write <= x"C8480000";
end if;
if first_state_sram_input_id = 9079 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 9080 then
	sram_write <= x"C8460004";
end if;
if first_state_sram_input_id = 9081 then
	sram_write <= x"C8680004";
end if;
if first_state_sram_input_id = 9082 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 9083 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 9084 then
	sram_write <= x"C8460008";
end if;
if first_state_sram_input_id = 9085 then
	sram_write <= x"C8680008";
end if;
if first_state_sram_input_id = 9086 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 9087 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 9088 then
	sram_write <= x"8E208E54";
end if;
if first_state_sram_input_id = 9089 then
	sram_write <= x"C8400018";
end if;
if first_state_sram_input_id = 9090 then
	sram_write <= x"C45C0078";
end if;
if first_state_sram_input_id = 9091 then
	sram_write <= x"CC3C0080";
end if;
if first_state_sram_input_id = 9092 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 9093 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 9094 then
	sram_write <= x"03DC0090";
end if;
if first_state_sram_input_id = 9095 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 9096 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 9097 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 9098 then
	sram_write <= x"07DC0090";
end if;
if first_state_sram_input_id = 9099 then
	sram_write <= x"C85C0080";
end if;
if first_state_sram_input_id = 9100 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 9101 then
	sram_write <= x"C03C0078";
end if;
if first_state_sram_input_id = 9102 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 9103 then
	sram_write <= x"03DC0090";
end if;
if first_state_sram_input_id = 9104 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 9105 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 9106 then
	sram_write <= x"82008034";
end if;
if first_state_sram_input_id = 9107 then
	sram_write <= x"07DC0090";
end if;
if first_state_sram_input_id = 9108 then
	sram_write <= x"82008EA4";
end if;
if first_state_sram_input_id = 9109 then
	sram_write <= x"C04201DC";
end if;
if first_state_sram_input_id = 9110 then
	sram_write <= x"C8400014";
end if;
if first_state_sram_input_id = 9111 then
	sram_write <= x"C45C0088";
end if;
if first_state_sram_input_id = 9112 then
	sram_write <= x"CC3C0080";
end if;
if first_state_sram_input_id = 9113 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 9114 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 9115 then
	sram_write <= x"03DC0094";
end if;
if first_state_sram_input_id = 9116 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 9117 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 9118 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 9119 then
	sram_write <= x"07DC0094";
end if;
if first_state_sram_input_id = 9120 then
	sram_write <= x"C85C0080";
end if;
if first_state_sram_input_id = 9121 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 9122 then
	sram_write <= x"C03C0088";
end if;
if first_state_sram_input_id = 9123 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 9124 then
	sram_write <= x"03DC0094";
end if;
if first_state_sram_input_id = 9125 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 9126 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 9127 then
	sram_write <= x"82008034";
end if;
if first_state_sram_input_id = 9128 then
	sram_write <= x"07DC0094";
end if;
if first_state_sram_input_id = 9129 then
	sram_write <= x"02800074";
end if;
if first_state_sram_input_id = 9130 then
	sram_write <= x"C03C0074";
end if;
if first_state_sram_input_id = 9131 then
	sram_write <= x"C05C000C";
end if;
if first_state_sram_input_id = 9132 then
	sram_write <= x"C07C0010";
end if;
if first_state_sram_input_id = 9133 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 9134 then
	sram_write <= x"03DC0094";
end if;
if first_state_sram_input_id = 9135 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 9136 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 9137 then
	sram_write <= x"82008280";
end if;
if first_state_sram_input_id = 9138 then
	sram_write <= x"07DC0094";
end if;
if first_state_sram_input_id = 9139 then
	sram_write <= x"82008ED0";
end if;
if first_state_sram_input_id = 9140 then
	sram_write <= x"022002EC";
end if;
if first_state_sram_input_id = 9141 then
	sram_write <= x"C05C0008";
end if;
if first_state_sram_input_id = 9142 then
	sram_write <= x"22440220";
end if;
if first_state_sram_input_id = 9143 then
	sram_write <= x"C07C0004";
end if;
if first_state_sram_input_id = 9144 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 9145 then
	sram_write <= x"C8220000";
end if;
if first_state_sram_input_id = 9146 then
	sram_write <= x"C8440000";
end if;
if first_state_sram_input_id = 9147 then
	sram_write <= x"C07C0000";
end if;
if first_state_sram_input_id = 9148 then
	sram_write <= x"C8660000";
end if;
if first_state_sram_input_id = 9149 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 9150 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 9151 then
	sram_write <= x"CC220000";
end if;
if first_state_sram_input_id = 9152 then
	sram_write <= x"C8220004";
end if;
if first_state_sram_input_id = 9153 then
	sram_write <= x"C8440004";
end if;
if first_state_sram_input_id = 9154 then
	sram_write <= x"C8660004";
end if;
if first_state_sram_input_id = 9155 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 9156 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 9157 then
	sram_write <= x"CC220004";
end if;
if first_state_sram_input_id = 9158 then
	sram_write <= x"C8220008";
end if;
if first_state_sram_input_id = 9159 then
	sram_write <= x"C8440008";
end if;
if first_state_sram_input_id = 9160 then
	sram_write <= x"C8660008";
end if;
if first_state_sram_input_id = 9161 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 9162 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 9163 then
	sram_write <= x"CC220008";
end if;
if first_state_sram_input_id = 9164 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 9165 then
	sram_write <= x"22C20220";
end if;
if first_state_sram_input_id = 9166 then
	sram_write <= x"D044C000";
end if;
if first_state_sram_input_id = 9167 then
	sram_write <= x"C0440014";
end if;
if first_state_sram_input_id = 9168 then
	sram_write <= x"06C20001";
end if;
if first_state_sram_input_id = 9169 then
	sram_write <= x"22CC0220";
end if;
if first_state_sram_input_id = 9170 then
	sram_write <= x"D0C6C000";
end if;
if first_state_sram_input_id = 9171 then
	sram_write <= x"C0CC0014";
end if;
if first_state_sram_input_id = 9172 then
	sram_write <= x"22E20220";
end if;
if first_state_sram_input_id = 9173 then
	sram_write <= x"D0E6E000";
end if;
if first_state_sram_input_id = 9174 then
	sram_write <= x"C0EE0014";
end if;
if first_state_sram_input_id = 9175 then
	sram_write <= x"03020001";
end if;
if first_state_sram_input_id = 9176 then
	sram_write <= x"23100220";
end if;
if first_state_sram_input_id = 9177 then
	sram_write <= x"D1070000";
end if;
if first_state_sram_input_id = 9178 then
	sram_write <= x"C1100014";
end if;
if first_state_sram_input_id = 9179 then
	sram_write <= x"23220220";
end if;
if first_state_sram_input_id = 9180 then
	sram_write <= x"D0892000";
end if;
if first_state_sram_input_id = 9181 then
	sram_write <= x"C0880014";
end if;
if first_state_sram_input_id = 9182 then
	sram_write <= x"032002E0";
end if;
if first_state_sram_input_id = 9183 then
	sram_write <= x"234A0220";
end if;
if first_state_sram_input_id = 9184 then
	sram_write <= x"D0454000";
end if;
if first_state_sram_input_id = 9185 then
	sram_write <= x"C8240000";
end if;
if first_state_sram_input_id = 9186 then
	sram_write <= x"CC320000";
end if;
if first_state_sram_input_id = 9187 then
	sram_write <= x"C8240004";
end if;
if first_state_sram_input_id = 9188 then
	sram_write <= x"CC320004";
end if;
if first_state_sram_input_id = 9189 then
	sram_write <= x"C8240008";
end if;
if first_state_sram_input_id = 9190 then
	sram_write <= x"CC320008";
end if;
if first_state_sram_input_id = 9191 then
	sram_write <= x"224A0220";
end if;
if first_state_sram_input_id = 9192 then
	sram_write <= x"D04C4000";
end if;
if first_state_sram_input_id = 9193 then
	sram_write <= x"C8320000";
end if;
if first_state_sram_input_id = 9194 then
	sram_write <= x"C8440000";
end if;
if first_state_sram_input_id = 9195 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 9196 then
	sram_write <= x"CC320000";
end if;
if first_state_sram_input_id = 9197 then
	sram_write <= x"C8320004";
end if;
if first_state_sram_input_id = 9198 then
	sram_write <= x"C8440004";
end if;
if first_state_sram_input_id = 9199 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 9200 then
	sram_write <= x"CC320004";
end if;
if first_state_sram_input_id = 9201 then
	sram_write <= x"C8320008";
end if;
if first_state_sram_input_id = 9202 then
	sram_write <= x"C8440008";
end if;
if first_state_sram_input_id = 9203 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 9204 then
	sram_write <= x"CC320008";
end if;
if first_state_sram_input_id = 9205 then
	sram_write <= x"224A0220";
end if;
if first_state_sram_input_id = 9206 then
	sram_write <= x"D04E4000";
end if;
if first_state_sram_input_id = 9207 then
	sram_write <= x"C8320000";
end if;
if first_state_sram_input_id = 9208 then
	sram_write <= x"C8440000";
end if;
if first_state_sram_input_id = 9209 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 9210 then
	sram_write <= x"CC320000";
end if;
if first_state_sram_input_id = 9211 then
	sram_write <= x"C8320004";
end if;
if first_state_sram_input_id = 9212 then
	sram_write <= x"C8440004";
end if;
if first_state_sram_input_id = 9213 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 9214 then
	sram_write <= x"CC320004";
end if;
if first_state_sram_input_id = 9215 then
	sram_write <= x"C8320008";
end if;
if first_state_sram_input_id = 9216 then
	sram_write <= x"C8440008";
end if;
if first_state_sram_input_id = 9217 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 9218 then
	sram_write <= x"CC320008";
end if;
if first_state_sram_input_id = 9219 then
	sram_write <= x"224A0220";
end if;
if first_state_sram_input_id = 9220 then
	sram_write <= x"D0504000";
end if;
if first_state_sram_input_id = 9221 then
	sram_write <= x"C8320000";
end if;
if first_state_sram_input_id = 9222 then
	sram_write <= x"C8440000";
end if;
if first_state_sram_input_id = 9223 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 9224 then
	sram_write <= x"CC320000";
end if;
if first_state_sram_input_id = 9225 then
	sram_write <= x"C8320004";
end if;
if first_state_sram_input_id = 9226 then
	sram_write <= x"C8440004";
end if;
if first_state_sram_input_id = 9227 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 9228 then
	sram_write <= x"CC320004";
end if;
if first_state_sram_input_id = 9229 then
	sram_write <= x"C8320008";
end if;
if first_state_sram_input_id = 9230 then
	sram_write <= x"C8440008";
end if;
if first_state_sram_input_id = 9231 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 9232 then
	sram_write <= x"CC320008";
end if;
if first_state_sram_input_id = 9233 then
	sram_write <= x"224A0220";
end if;
if first_state_sram_input_id = 9234 then
	sram_write <= x"D0484000";
end if;
if first_state_sram_input_id = 9235 then
	sram_write <= x"C8320000";
end if;
if first_state_sram_input_id = 9236 then
	sram_write <= x"C8440000";
end if;
if first_state_sram_input_id = 9237 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 9238 then
	sram_write <= x"CC320000";
end if;
if first_state_sram_input_id = 9239 then
	sram_write <= x"C8320004";
end if;
if first_state_sram_input_id = 9240 then
	sram_write <= x"C8440004";
end if;
if first_state_sram_input_id = 9241 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 9242 then
	sram_write <= x"CC320004";
end if;
if first_state_sram_input_id = 9243 then
	sram_write <= x"C8320008";
end if;
if first_state_sram_input_id = 9244 then
	sram_write <= x"C8440008";
end if;
if first_state_sram_input_id = 9245 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 9246 then
	sram_write <= x"CC320008";
end if;
if first_state_sram_input_id = 9247 then
	sram_write <= x"22220220";
end if;
if first_state_sram_input_id = 9248 then
	sram_write <= x"D0262000";
end if;
if first_state_sram_input_id = 9249 then
	sram_write <= x"C0220010";
end if;
if first_state_sram_input_id = 9250 then
	sram_write <= x"024002EC";
end if;
if first_state_sram_input_id = 9251 then
	sram_write <= x"226A0220";
end if;
if first_state_sram_input_id = 9252 then
	sram_write <= x"D0226000";
end if;
if first_state_sram_input_id = 9253 then
	sram_write <= x"C8240000";
end if;
if first_state_sram_input_id = 9254 then
	sram_write <= x"C8420000";
end if;
if first_state_sram_input_id = 9255 then
	sram_write <= x"C8720000";
end if;
if first_state_sram_input_id = 9256 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 9257 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 9258 then
	sram_write <= x"CC240000";
end if;
if first_state_sram_input_id = 9259 then
	sram_write <= x"C8240004";
end if;
if first_state_sram_input_id = 9260 then
	sram_write <= x"C8420004";
end if;
if first_state_sram_input_id = 9261 then
	sram_write <= x"C8720004";
end if;
if first_state_sram_input_id = 9262 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 9263 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 9264 then
	sram_write <= x"CC240004";
end if;
if first_state_sram_input_id = 9265 then
	sram_write <= x"C8240008";
end if;
if first_state_sram_input_id = 9266 then
	sram_write <= x"C8420008";
end if;
if first_state_sram_input_id = 9267 then
	sram_write <= x"C8720008";
end if;
if first_state_sram_input_id = 9268 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 9269 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 9270 then
	sram_write <= x"CC240008";
end if;
if first_state_sram_input_id = 9271 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 9272 then
	sram_write <= x"02600004";
end if;
if first_state_sram_input_id = 9273 then
	sram_write <= x"86649258";
end if;
if first_state_sram_input_id = 9274 then
	sram_write <= x"C0620008";
end if;
if first_state_sram_input_id = 9275 then
	sram_write <= x"22840220";
end if;
if first_state_sram_input_id = 9276 then
	sram_write <= x"D0668000";
end if;
if first_state_sram_input_id = 9277 then
	sram_write <= x"86609254";
end if;
if first_state_sram_input_id = 9278 then
	sram_write <= x"C062000C";
end if;
if first_state_sram_input_id = 9279 then
	sram_write <= x"22840220";
end if;
if first_state_sram_input_id = 9280 then
	sram_write <= x"D0668000";
end if;
if first_state_sram_input_id = 9281 then
	sram_write <= x"C43C0000";
end if;
if first_state_sram_input_id = 9282 then
	sram_write <= x"826091EC";
end if;
if first_state_sram_input_id = 9283 then
	sram_write <= x"C0620014";
end if;
if first_state_sram_input_id = 9284 then
	sram_write <= x"C082001C";
end if;
if first_state_sram_input_id = 9285 then
	sram_write <= x"C0A20004";
end if;
if first_state_sram_input_id = 9286 then
	sram_write <= x"C0C20010";
end if;
if first_state_sram_input_id = 9287 then
	sram_write <= x"02E002E0";
end if;
if first_state_sram_input_id = 9288 then
	sram_write <= x"23040220";
end if;
if first_state_sram_input_id = 9289 then
	sram_write <= x"D0670000";
end if;
if first_state_sram_input_id = 9290 then
	sram_write <= x"C8260000";
end if;
if first_state_sram_input_id = 9291 then
	sram_write <= x"CC2E0000";
end if;
if first_state_sram_input_id = 9292 then
	sram_write <= x"C8260004";
end if;
if first_state_sram_input_id = 9293 then
	sram_write <= x"CC2E0004";
end if;
if first_state_sram_input_id = 9294 then
	sram_write <= x"C8260008";
end if;
if first_state_sram_input_id = 9295 then
	sram_write <= x"CC2E0008";
end if;
if first_state_sram_input_id = 9296 then
	sram_write <= x"C0620018";
end if;
if first_state_sram_input_id = 9297 then
	sram_write <= x"C0660000";
end if;
if first_state_sram_input_id = 9298 then
	sram_write <= x"23040220";
end if;
if first_state_sram_input_id = 9299 then
	sram_write <= x"D0890000";
end if;
if first_state_sram_input_id = 9300 then
	sram_write <= x"23040220";
end if;
if first_state_sram_input_id = 9301 then
	sram_write <= x"D0AB0000";
end if;
if first_state_sram_input_id = 9302 then
	sram_write <= x"C4FC0004";
end if;
if first_state_sram_input_id = 9303 then
	sram_write <= x"C4DC0008";
end if;
if first_state_sram_input_id = 9304 then
	sram_write <= x"C45C000C";
end if;
if first_state_sram_input_id = 9305 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 9306 then
	sram_write <= x"00480000";
end if;
if first_state_sram_input_id = 9307 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 9308 then
	sram_write <= x"006A0000";
end if;
if first_state_sram_input_id = 9309 then
	sram_write <= x"03DC0018";
end if;
if first_state_sram_input_id = 9310 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 9311 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 9312 then
	sram_write <= x"82008494";
end if;
if first_state_sram_input_id = 9313 then
	sram_write <= x"07DC0018";
end if;
if first_state_sram_input_id = 9314 then
	sram_write <= x"022002EC";
end if;
if first_state_sram_input_id = 9315 then
	sram_write <= x"C05C000C";
end if;
if first_state_sram_input_id = 9316 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 9317 then
	sram_write <= x"C09C0008";
end if;
if first_state_sram_input_id = 9318 then
	sram_write <= x"D0686000";
end if;
if first_state_sram_input_id = 9319 then
	sram_write <= x"C8220000";
end if;
if first_state_sram_input_id = 9320 then
	sram_write <= x"C8460000";
end if;
if first_state_sram_input_id = 9321 then
	sram_write <= x"C09C0004";
end if;
if first_state_sram_input_id = 9322 then
	sram_write <= x"C8680000";
end if;
if first_state_sram_input_id = 9323 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 9324 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 9325 then
	sram_write <= x"CC220000";
end if;
if first_state_sram_input_id = 9326 then
	sram_write <= x"C8220004";
end if;
if first_state_sram_input_id = 9327 then
	sram_write <= x"C8460004";
end if;
if first_state_sram_input_id = 9328 then
	sram_write <= x"C8680004";
end if;
if first_state_sram_input_id = 9329 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 9330 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 9331 then
	sram_write <= x"CC220004";
end if;
if first_state_sram_input_id = 9332 then
	sram_write <= x"C8220008";
end if;
if first_state_sram_input_id = 9333 then
	sram_write <= x"C8460008";
end if;
if first_state_sram_input_id = 9334 then
	sram_write <= x"C8680008";
end if;
if first_state_sram_input_id = 9335 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 9336 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 9337 then
	sram_write <= x"CC220008";
end if;
if first_state_sram_input_id = 9338 then
	sram_write <= x"820091EC";
end if;
if first_state_sram_input_id = 9339 then
	sram_write <= x"02440001";
end if;
if first_state_sram_input_id = 9340 then
	sram_write <= x"02200004";
end if;
if first_state_sram_input_id = 9341 then
	sram_write <= x"86249250";
end if;
if first_state_sram_input_id = 9342 then
	sram_write <= x"C03C0000";
end if;
if first_state_sram_input_id = 9343 then
	sram_write <= x"C0620008";
end if;
if first_state_sram_input_id = 9344 then
	sram_write <= x"22840220";
end if;
if first_state_sram_input_id = 9345 then
	sram_write <= x"D0668000";
end if;
if first_state_sram_input_id = 9346 then
	sram_write <= x"8660924C";
end if;
if first_state_sram_input_id = 9347 then
	sram_write <= x"C062000C";
end if;
if first_state_sram_input_id = 9348 then
	sram_write <= x"22840220";
end if;
if first_state_sram_input_id = 9349 then
	sram_write <= x"D0668000";
end if;
if first_state_sram_input_id = 9350 then
	sram_write <= x"C45C0010";
end if;
if first_state_sram_input_id = 9351 then
	sram_write <= x"8260923C";
end if;
if first_state_sram_input_id = 9352 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 9353 then
	sram_write <= x"03DC001C";
end if;
if first_state_sram_input_id = 9354 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 9355 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 9356 then
	sram_write <= x"8200874C";
end if;
if first_state_sram_input_id = 9357 then
	sram_write <= x"07DC001C";
end if;
if first_state_sram_input_id = 9358 then
	sram_write <= x"8200923C";
end if;
if first_state_sram_input_id = 9359 then
	sram_write <= x"C03C0010";
end if;
if first_state_sram_input_id = 9360 then
	sram_write <= x"02420001";
end if;
if first_state_sram_input_id = 9361 then
	sram_write <= x"C03C0000";
end if;
if first_state_sram_input_id = 9362 then
	sram_write <= x"820090E0";
end if;
if first_state_sram_input_id = 9363 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 9364 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 9365 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 9366 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 9367 then
	sram_write <= x"22E20220";
end if;
if first_state_sram_input_id = 9368 then
	sram_write <= x"D0E8E000";
end if;
if first_state_sram_input_id = 9369 then
	sram_write <= x"03000004";
end if;
if first_state_sram_input_id = 9370 then
	sram_write <= x"870C9528";
end if;
if first_state_sram_input_id = 9371 then
	sram_write <= x"C10E0008";
end if;
if first_state_sram_input_id = 9372 then
	sram_write <= x"232C0220";
end if;
if first_state_sram_input_id = 9373 then
	sram_write <= x"D1112000";
end if;
if first_state_sram_input_id = 9374 then
	sram_write <= x"87009524";
end if;
if first_state_sram_input_id = 9375 then
	sram_write <= x"C10E0008";
end if;
if first_state_sram_input_id = 9376 then
	sram_write <= x"232C0220";
end if;
if first_state_sram_input_id = 9377 then
	sram_write <= x"D1112000";
end if;
if first_state_sram_input_id = 9378 then
	sram_write <= x"23220220";
end if;
if first_state_sram_input_id = 9379 then
	sram_write <= x"D1272000";
end if;
if first_state_sram_input_id = 9380 then
	sram_write <= x"C1320008";
end if;
if first_state_sram_input_id = 9381 then
	sram_write <= x"234C0220";
end if;
if first_state_sram_input_id = 9382 then
	sram_write <= x"D1334000";
end if;
if first_state_sram_input_id = 9383 then
	sram_write <= x"833092A8";
end if;
if first_state_sram_input_id = 9384 then
	sram_write <= x"03000000";
end if;
if first_state_sram_input_id = 9385 then
	sram_write <= x"82009314";
end if;
if first_state_sram_input_id = 9386 then
	sram_write <= x"23220220";
end if;
if first_state_sram_input_id = 9387 then
	sram_write <= x"D12B2000";
end if;
if first_state_sram_input_id = 9388 then
	sram_write <= x"C1320008";
end if;
if first_state_sram_input_id = 9389 then
	sram_write <= x"234C0220";
end if;
if first_state_sram_input_id = 9390 then
	sram_write <= x"D1334000";
end if;
if first_state_sram_input_id = 9391 then
	sram_write <= x"833092C8";
end if;
if first_state_sram_input_id = 9392 then
	sram_write <= x"03000000";
end if;
if first_state_sram_input_id = 9393 then
	sram_write <= x"82009314";
end if;
if first_state_sram_input_id = 9394 then
	sram_write <= x"07220001";
end if;
if first_state_sram_input_id = 9395 then
	sram_write <= x"23320220";
end if;
if first_state_sram_input_id = 9396 then
	sram_write <= x"D1292000";
end if;
if first_state_sram_input_id = 9397 then
	sram_write <= x"C1320008";
end if;
if first_state_sram_input_id = 9398 then
	sram_write <= x"234C0220";
end if;
if first_state_sram_input_id = 9399 then
	sram_write <= x"D1334000";
end if;
if first_state_sram_input_id = 9400 then
	sram_write <= x"833092EC";
end if;
if first_state_sram_input_id = 9401 then
	sram_write <= x"03000000";
end if;
if first_state_sram_input_id = 9402 then
	sram_write <= x"82009314";
end if;
if first_state_sram_input_id = 9403 then
	sram_write <= x"03220001";
end if;
if first_state_sram_input_id = 9404 then
	sram_write <= x"23320220";
end if;
if first_state_sram_input_id = 9405 then
	sram_write <= x"D1292000";
end if;
if first_state_sram_input_id = 9406 then
	sram_write <= x"C1320008";
end if;
if first_state_sram_input_id = 9407 then
	sram_write <= x"234C0220";
end if;
if first_state_sram_input_id = 9408 then
	sram_write <= x"D1334000";
end if;
if first_state_sram_input_id = 9409 then
	sram_write <= x"83309310";
end if;
if first_state_sram_input_id = 9410 then
	sram_write <= x"03000000";
end if;
if first_state_sram_input_id = 9411 then
	sram_write <= x"82009314";
end if;
if first_state_sram_input_id = 9412 then
	sram_write <= x"03000001";
end if;
if first_state_sram_input_id = 9413 then
	sram_write <= x"830094B8";
end if;
if first_state_sram_input_id = 9414 then
	sram_write <= x"C0EE000C";
end if;
if first_state_sram_input_id = 9415 then
	sram_write <= x"230C0220";
end if;
if first_state_sram_input_id = 9416 then
	sram_write <= x"D0EF0000";
end if;
if first_state_sram_input_id = 9417 then
	sram_write <= x"C45C0000";
end if;
if first_state_sram_input_id = 9418 then
	sram_write <= x"C4BC0004";
end if;
if first_state_sram_input_id = 9419 then
	sram_write <= x"C47C0008";
end if;
if first_state_sram_input_id = 9420 then
	sram_write <= x"C49C000C";
end if;
if first_state_sram_input_id = 9421 then
	sram_write <= x"C43C0010";
end if;
if first_state_sram_input_id = 9422 then
	sram_write <= x"C4DC0014";
end if;
if first_state_sram_input_id = 9423 then
	sram_write <= x"82E0936C";
end if;
if first_state_sram_input_id = 9424 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 9425 then
	sram_write <= x"00460000";
end if;
if first_state_sram_input_id = 9426 then
	sram_write <= x"00680000";
end if;
if first_state_sram_input_id = 9427 then
	sram_write <= x"008A0000";
end if;
if first_state_sram_input_id = 9428 then
	sram_write <= x"00AC0000";
end if;
if first_state_sram_input_id = 9429 then
	sram_write <= x"03DC0020";
end if;
if first_state_sram_input_id = 9430 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 9431 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 9432 then
	sram_write <= x"82008F34";
end if;
if first_state_sram_input_id = 9433 then
	sram_write <= x"07DC0020";
end if;
if first_state_sram_input_id = 9434 then
	sram_write <= x"8200936C";
end if;
if first_state_sram_input_id = 9435 then
	sram_write <= x"C03C0014";
end if;
if first_state_sram_input_id = 9436 then
	sram_write <= x"02420001";
end if;
if first_state_sram_input_id = 9437 then
	sram_write <= x"C03C0010";
end if;
if first_state_sram_input_id = 9438 then
	sram_write <= x"22620220";
end if;
if first_state_sram_input_id = 9439 then
	sram_write <= x"C09C000C";
end if;
if first_state_sram_input_id = 9440 then
	sram_write <= x"D0686000";
end if;
if first_state_sram_input_id = 9441 then
	sram_write <= x"02A00004";
end if;
if first_state_sram_input_id = 9442 then
	sram_write <= x"86A494B4";
end if;
if first_state_sram_input_id = 9443 then
	sram_write <= x"C0A60008";
end if;
if first_state_sram_input_id = 9444 then
	sram_write <= x"22C40220";
end if;
if first_state_sram_input_id = 9445 then
	sram_write <= x"D0AAC000";
end if;
if first_state_sram_input_id = 9446 then
	sram_write <= x"86A094B0";
end if;
if first_state_sram_input_id = 9447 then
	sram_write <= x"C0A60008";
end if;
if first_state_sram_input_id = 9448 then
	sram_write <= x"22C40220";
end if;
if first_state_sram_input_id = 9449 then
	sram_write <= x"D0AAC000";
end if;
if first_state_sram_input_id = 9450 then
	sram_write <= x"22C20220";
end if;
if first_state_sram_input_id = 9451 then
	sram_write <= x"C0FC0008";
end if;
if first_state_sram_input_id = 9452 then
	sram_write <= x"D0CEC000";
end if;
if first_state_sram_input_id = 9453 then
	sram_write <= x"C0CC0008";
end if;
if first_state_sram_input_id = 9454 then
	sram_write <= x"23040220";
end if;
if first_state_sram_input_id = 9455 then
	sram_write <= x"D0CD0000";
end if;
if first_state_sram_input_id = 9456 then
	sram_write <= x"82CA93CC";
end if;
if first_state_sram_input_id = 9457 then
	sram_write <= x"02A00000";
end if;
if first_state_sram_input_id = 9458 then
	sram_write <= x"8200943C";
end if;
if first_state_sram_input_id = 9459 then
	sram_write <= x"22C20220";
end if;
if first_state_sram_input_id = 9460 then
	sram_write <= x"C11C0004";
end if;
if first_state_sram_input_id = 9461 then
	sram_write <= x"D0D0C000";
end if;
if first_state_sram_input_id = 9462 then
	sram_write <= x"C0CC0008";
end if;
if first_state_sram_input_id = 9463 then
	sram_write <= x"23240220";
end if;
if first_state_sram_input_id = 9464 then
	sram_write <= x"D0CD2000";
end if;
if first_state_sram_input_id = 9465 then
	sram_write <= x"82CA93F0";
end if;
if first_state_sram_input_id = 9466 then
	sram_write <= x"02A00000";
end if;
if first_state_sram_input_id = 9467 then
	sram_write <= x"8200943C";
end if;
if first_state_sram_input_id = 9468 then
	sram_write <= x"06C20001";
end if;
if first_state_sram_input_id = 9469 then
	sram_write <= x"22CC0220";
end if;
if first_state_sram_input_id = 9470 then
	sram_write <= x"D0C8C000";
end if;
if first_state_sram_input_id = 9471 then
	sram_write <= x"C0CC0008";
end if;
if first_state_sram_input_id = 9472 then
	sram_write <= x"23240220";
end if;
if first_state_sram_input_id = 9473 then
	sram_write <= x"D0CD2000";
end if;
if first_state_sram_input_id = 9474 then
	sram_write <= x"82CA9414";
end if;
if first_state_sram_input_id = 9475 then
	sram_write <= x"02A00000";
end if;
if first_state_sram_input_id = 9476 then
	sram_write <= x"8200943C";
end if;
if first_state_sram_input_id = 9477 then
	sram_write <= x"02C20001";
end if;
if first_state_sram_input_id = 9478 then
	sram_write <= x"22CC0220";
end if;
if first_state_sram_input_id = 9479 then
	sram_write <= x"D0C8C000";
end if;
if first_state_sram_input_id = 9480 then
	sram_write <= x"C0CC0008";
end if;
if first_state_sram_input_id = 9481 then
	sram_write <= x"23240220";
end if;
if first_state_sram_input_id = 9482 then
	sram_write <= x"D0CD2000";
end if;
if first_state_sram_input_id = 9483 then
	sram_write <= x"82CA9438";
end if;
if first_state_sram_input_id = 9484 then
	sram_write <= x"02A00000";
end if;
if first_state_sram_input_id = 9485 then
	sram_write <= x"8200943C";
end if;
if first_state_sram_input_id = 9486 then
	sram_write <= x"02A00001";
end if;
if first_state_sram_input_id = 9487 then
	sram_write <= x"82A094A8";
end if;
if first_state_sram_input_id = 9488 then
	sram_write <= x"C066000C";
end if;
if first_state_sram_input_id = 9489 then
	sram_write <= x"22A40220";
end if;
if first_state_sram_input_id = 9490 then
	sram_write <= x"D066A000";
end if;
if first_state_sram_input_id = 9491 then
	sram_write <= x"C45C0018";
end if;
if first_state_sram_input_id = 9492 then
	sram_write <= x"82609488";
end if;
if first_state_sram_input_id = 9493 then
	sram_write <= x"C07C0004";
end if;
if first_state_sram_input_id = 9494 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 9495 then
	sram_write <= x"00A40000";
end if;
if first_state_sram_input_id = 9496 then
	sram_write <= x"004E0000";
end if;
if first_state_sram_input_id = 9497 then
	sram_write <= x"01280000";
end if;
if first_state_sram_input_id = 9498 then
	sram_write <= x"00860000";
end if;
if first_state_sram_input_id = 9499 then
	sram_write <= x"00720000";
end if;
if first_state_sram_input_id = 9500 then
	sram_write <= x"03DC0024";
end if;
if first_state_sram_input_id = 9501 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 9502 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 9503 then
	sram_write <= x"82008F34";
end if;
if first_state_sram_input_id = 9504 then
	sram_write <= x"07DC0024";
end if;
if first_state_sram_input_id = 9505 then
	sram_write <= x"82009488";
end if;
if first_state_sram_input_id = 9506 then
	sram_write <= x"C03C0018";
end if;
if first_state_sram_input_id = 9507 then
	sram_write <= x"02C20001";
end if;
if first_state_sram_input_id = 9508 then
	sram_write <= x"C03C0010";
end if;
if first_state_sram_input_id = 9509 then
	sram_write <= x"C05C0000";
end if;
if first_state_sram_input_id = 9510 then
	sram_write <= x"C07C0008";
end if;
if first_state_sram_input_id = 9511 then
	sram_write <= x"C09C000C";
end if;
if first_state_sram_input_id = 9512 then
	sram_write <= x"C0BC0004";
end if;
if first_state_sram_input_id = 9513 then
	sram_write <= x"8200925C";
end if;
if first_state_sram_input_id = 9514 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 9515 then
	sram_write <= x"820090E0";
end if;
if first_state_sram_input_id = 9516 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 9517 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 9518 then
	sram_write <= x"02200004";
end if;
if first_state_sram_input_id = 9519 then
	sram_write <= x"862C9520";
end if;
if first_state_sram_input_id = 9520 then
	sram_write <= x"C02E0008";
end if;
if first_state_sram_input_id = 9521 then
	sram_write <= x"224C0220";
end if;
if first_state_sram_input_id = 9522 then
	sram_write <= x"D0224000";
end if;
if first_state_sram_input_id = 9523 then
	sram_write <= x"8620951C";
end if;
if first_state_sram_input_id = 9524 then
	sram_write <= x"C02E000C";
end if;
if first_state_sram_input_id = 9525 then
	sram_write <= x"224C0220";
end if;
if first_state_sram_input_id = 9526 then
	sram_write <= x"D0224000";
end if;
if first_state_sram_input_id = 9527 then
	sram_write <= x"C4FC001C";
end if;
if first_state_sram_input_id = 9528 then
	sram_write <= x"C4DC0014";
end if;
if first_state_sram_input_id = 9529 then
	sram_write <= x"8220950C";
end if;
if first_state_sram_input_id = 9530 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 9531 then
	sram_write <= x"004C0000";
end if;
if first_state_sram_input_id = 9532 then
	sram_write <= x"002E0000";
end if;
if first_state_sram_input_id = 9533 then
	sram_write <= x"03DC0028";
end if;
if first_state_sram_input_id = 9534 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 9535 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 9536 then
	sram_write <= x"8200874C";
end if;
if first_state_sram_input_id = 9537 then
	sram_write <= x"07DC0028";
end if;
if first_state_sram_input_id = 9538 then
	sram_write <= x"8200950C";
end if;
if first_state_sram_input_id = 9539 then
	sram_write <= x"C03C0014";
end if;
if first_state_sram_input_id = 9540 then
	sram_write <= x"02420001";
end if;
if first_state_sram_input_id = 9541 then
	sram_write <= x"C03C001C";
end if;
if first_state_sram_input_id = 9542 then
	sram_write <= x"820090E0";
end if;
if first_state_sram_input_id = 9543 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 9544 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 9545 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 9546 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 9547 then
	sram_write <= x"02600004";
end if;
if first_state_sram_input_id = 9548 then
	sram_write <= x"8664986C";
end if;
if first_state_sram_input_id = 9549 then
	sram_write <= x"C0620008";
end if;
if first_state_sram_input_id = 9550 then
	sram_write <= x"22840220";
end if;
if first_state_sram_input_id = 9551 then
	sram_write <= x"D0668000";
end if;
if first_state_sram_input_id = 9552 then
	sram_write <= x"86609868";
end if;
if first_state_sram_input_id = 9553 then
	sram_write <= x"C062000C";
end if;
if first_state_sram_input_id = 9554 then
	sram_write <= x"22840220";
end if;
if first_state_sram_input_id = 9555 then
	sram_write <= x"D0668000";
end if;
if first_state_sram_input_id = 9556 then
	sram_write <= x"C45C0000";
end if;
if first_state_sram_input_id = 9557 then
	sram_write <= x"8260964C";
end if;
if first_state_sram_input_id = 9558 then
	sram_write <= x"C0620018";
end if;
if first_state_sram_input_id = 9559 then
	sram_write <= x"C0660000";
end if;
if first_state_sram_input_id = 9560 then
	sram_write <= x"028002E0";
end if;
if first_state_sram_input_id = 9561 then
	sram_write <= x"CC080000";
end if;
if first_state_sram_input_id = 9562 then
	sram_write <= x"CC080004";
end if;
if first_state_sram_input_id = 9563 then
	sram_write <= x"CC080008";
end if;
if first_state_sram_input_id = 9564 then
	sram_write <= x"C0A2001C";
end if;
if first_state_sram_input_id = 9565 then
	sram_write <= x"C0C20004";
end if;
if first_state_sram_input_id = 9566 then
	sram_write <= x"02E00354";
end if;
if first_state_sram_input_id = 9567 then
	sram_write <= x"22660220";
end if;
if first_state_sram_input_id = 9568 then
	sram_write <= x"D06E6000";
end if;
if first_state_sram_input_id = 9569 then
	sram_write <= x"22E40220";
end if;
if first_state_sram_input_id = 9570 then
	sram_write <= x"D0AAE000";
end if;
if first_state_sram_input_id = 9571 then
	sram_write <= x"22E40220";
end if;
if first_state_sram_input_id = 9572 then
	sram_write <= x"D0CCE000";
end if;
if first_state_sram_input_id = 9573 then
	sram_write <= x"02E00318";
end if;
if first_state_sram_input_id = 9574 then
	sram_write <= x"C82C0000";
end if;
if first_state_sram_input_id = 9575 then
	sram_write <= x"CC2E0000";
end if;
if first_state_sram_input_id = 9576 then
	sram_write <= x"C82C0004";
end if;
if first_state_sram_input_id = 9577 then
	sram_write <= x"CC2E0004";
end if;
if first_state_sram_input_id = 9578 then
	sram_write <= x"C82C0008";
end if;
if first_state_sram_input_id = 9579 then
	sram_write <= x"CC2E0008";
end if;
if first_state_sram_input_id = 9580 then
	sram_write <= x"02E000C4";
end if;
if first_state_sram_input_id = 9581 then
	sram_write <= x"C0EE0000";
end if;
if first_state_sram_input_id = 9582 then
	sram_write <= x"06EE0001";
end if;
if first_state_sram_input_id = 9583 then
	sram_write <= x"C49C0004";
end if;
if first_state_sram_input_id = 9584 then
	sram_write <= x"C43C0008";
end if;
if first_state_sram_input_id = 9585 then
	sram_write <= x"C4DC000C";
end if;
if first_state_sram_input_id = 9586 then
	sram_write <= x"C4BC0010";
end if;
if first_state_sram_input_id = 9587 then
	sram_write <= x"C47C0014";
end if;
if first_state_sram_input_id = 9588 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 9589 then
	sram_write <= x"004E0000";
end if;
if first_state_sram_input_id = 9590 then
	sram_write <= x"002C0000";
end if;
if first_state_sram_input_id = 9591 then
	sram_write <= x"03DC0020";
end if;
if first_state_sram_input_id = 9592 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 9593 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 9594 then
	sram_write <= x"8200462C";
end if;
if first_state_sram_input_id = 9595 then
	sram_write <= x"07DC0020";
end if;
if first_state_sram_input_id = 9596 then
	sram_write <= x"02800076";
end if;
if first_state_sram_input_id = 9597 then
	sram_write <= x"C03C0014";
end if;
if first_state_sram_input_id = 9598 then
	sram_write <= x"C05C0010";
end if;
if first_state_sram_input_id = 9599 then
	sram_write <= x"C07C000C";
end if;
if first_state_sram_input_id = 9600 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 9601 then
	sram_write <= x"03DC0020";
end if;
if first_state_sram_input_id = 9602 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 9603 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 9604 then
	sram_write <= x"82008280";
end if;
if first_state_sram_input_id = 9605 then
	sram_write <= x"07DC0020";
end if;
if first_state_sram_input_id = 9606 then
	sram_write <= x"C03C0008";
end if;
if first_state_sram_input_id = 9607 then
	sram_write <= x"C0420014";
end if;
if first_state_sram_input_id = 9608 then
	sram_write <= x"C07C0000";
end if;
if first_state_sram_input_id = 9609 then
	sram_write <= x"22860220";
end if;
if first_state_sram_input_id = 9610 then
	sram_write <= x"D0448000";
end if;
if first_state_sram_input_id = 9611 then
	sram_write <= x"C09C0004";
end if;
if first_state_sram_input_id = 9612 then
	sram_write <= x"C8280000";
end if;
if first_state_sram_input_id = 9613 then
	sram_write <= x"CC240000";
end if;
if first_state_sram_input_id = 9614 then
	sram_write <= x"C8280004";
end if;
if first_state_sram_input_id = 9615 then
	sram_write <= x"CC240004";
end if;
if first_state_sram_input_id = 9616 then
	sram_write <= x"C8280008";
end if;
if first_state_sram_input_id = 9617 then
	sram_write <= x"CC240008";
end if;
if first_state_sram_input_id = 9618 then
	sram_write <= x"8200964C";
end if;
if first_state_sram_input_id = 9619 then
	sram_write <= x"C05C0000";
end if;
if first_state_sram_input_id = 9620 then
	sram_write <= x"02440001";
end if;
if first_state_sram_input_id = 9621 then
	sram_write <= x"02600004";
end if;
if first_state_sram_input_id = 9622 then
	sram_write <= x"86649864";
end if;
if first_state_sram_input_id = 9623 then
	sram_write <= x"C0620008";
end if;
if first_state_sram_input_id = 9624 then
	sram_write <= x"22840220";
end if;
if first_state_sram_input_id = 9625 then
	sram_write <= x"D0668000";
end if;
if first_state_sram_input_id = 9626 then
	sram_write <= x"86609860";
end if;
if first_state_sram_input_id = 9627 then
	sram_write <= x"C062000C";
end if;
if first_state_sram_input_id = 9628 then
	sram_write <= x"22840220";
end if;
if first_state_sram_input_id = 9629 then
	sram_write <= x"D0668000";
end if;
if first_state_sram_input_id = 9630 then
	sram_write <= x"C45C0018";
end if;
if first_state_sram_input_id = 9631 then
	sram_write <= x"82609854";
end if;
if first_state_sram_input_id = 9632 then
	sram_write <= x"C0620018";
end if;
if first_state_sram_input_id = 9633 then
	sram_write <= x"C0660000";
end if;
if first_state_sram_input_id = 9634 then
	sram_write <= x"028002E0";
end if;
if first_state_sram_input_id = 9635 then
	sram_write <= x"CC080000";
end if;
if first_state_sram_input_id = 9636 then
	sram_write <= x"CC080004";
end if;
if first_state_sram_input_id = 9637 then
	sram_write <= x"CC080008";
end if;
if first_state_sram_input_id = 9638 then
	sram_write <= x"C0A2001C";
end if;
if first_state_sram_input_id = 9639 then
	sram_write <= x"C0C20004";
end if;
if first_state_sram_input_id = 9640 then
	sram_write <= x"02E00354";
end if;
if first_state_sram_input_id = 9641 then
	sram_write <= x"22660220";
end if;
if first_state_sram_input_id = 9642 then
	sram_write <= x"D06E6000";
end if;
if first_state_sram_input_id = 9643 then
	sram_write <= x"22E40220";
end if;
if first_state_sram_input_id = 9644 then
	sram_write <= x"D0AAE000";
end if;
if first_state_sram_input_id = 9645 then
	sram_write <= x"22E40220";
end if;
if first_state_sram_input_id = 9646 then
	sram_write <= x"D0CCE000";
end if;
if first_state_sram_input_id = 9647 then
	sram_write <= x"02E00318";
end if;
if first_state_sram_input_id = 9648 then
	sram_write <= x"C82C0000";
end if;
if first_state_sram_input_id = 9649 then
	sram_write <= x"CC2E0000";
end if;
if first_state_sram_input_id = 9650 then
	sram_write <= x"C82C0004";
end if;
if first_state_sram_input_id = 9651 then
	sram_write <= x"CC2E0004";
end if;
if first_state_sram_input_id = 9652 then
	sram_write <= x"C82C0008";
end if;
if first_state_sram_input_id = 9653 then
	sram_write <= x"CC2E0008";
end if;
if first_state_sram_input_id = 9654 then
	sram_write <= x"02E000C4";
end if;
if first_state_sram_input_id = 9655 then
	sram_write <= x"C0EE0000";
end if;
if first_state_sram_input_id = 9656 then
	sram_write <= x"06EE0001";
end if;
if first_state_sram_input_id = 9657 then
	sram_write <= x"C49C001C";
end if;
if first_state_sram_input_id = 9658 then
	sram_write <= x"C43C0008";
end if;
if first_state_sram_input_id = 9659 then
	sram_write <= x"C4DC0020";
end if;
if first_state_sram_input_id = 9660 then
	sram_write <= x"C4BC0024";
end if;
if first_state_sram_input_id = 9661 then
	sram_write <= x"C47C0028";
end if;
if first_state_sram_input_id = 9662 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 9663 then
	sram_write <= x"004E0000";
end if;
if first_state_sram_input_id = 9664 then
	sram_write <= x"002C0000";
end if;
if first_state_sram_input_id = 9665 then
	sram_write <= x"03DC0034";
end if;
if first_state_sram_input_id = 9666 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 9667 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 9668 then
	sram_write <= x"8200462C";
end if;
if first_state_sram_input_id = 9669 then
	sram_write <= x"07DC0034";
end if;
if first_state_sram_input_id = 9670 then
	sram_write <= x"C03C0028";
end if;
if first_state_sram_input_id = 9671 then
	sram_write <= x"C04201D8";
end if;
if first_state_sram_input_id = 9672 then
	sram_write <= x"C0640000";
end if;
if first_state_sram_input_id = 9673 then
	sram_write <= x"C8260000";
end if;
if first_state_sram_input_id = 9674 then
	sram_write <= x"C09C0024";
end if;
if first_state_sram_input_id = 9675 then
	sram_write <= x"C8480000";
end if;
if first_state_sram_input_id = 9676 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 9677 then
	sram_write <= x"C8460004";
end if;
if first_state_sram_input_id = 9678 then
	sram_write <= x"C8680004";
end if;
if first_state_sram_input_id = 9679 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 9680 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 9681 then
	sram_write <= x"C8460008";
end if;
if first_state_sram_input_id = 9682 then
	sram_write <= x"C8680008";
end if;
if first_state_sram_input_id = 9683 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 9684 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 9685 then
	sram_write <= x"8E2097A8";
end if;
if first_state_sram_input_id = 9686 then
	sram_write <= x"C8400018";
end if;
if first_state_sram_input_id = 9687 then
	sram_write <= x"C45C002C";
end if;
if first_state_sram_input_id = 9688 then
	sram_write <= x"CC3C0030";
end if;
if first_state_sram_input_id = 9689 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 9690 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 9691 then
	sram_write <= x"03DC0040";
end if;
if first_state_sram_input_id = 9692 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 9693 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 9694 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 9695 then
	sram_write <= x"07DC0040";
end if;
if first_state_sram_input_id = 9696 then
	sram_write <= x"C85C0030";
end if;
if first_state_sram_input_id = 9697 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 9698 then
	sram_write <= x"C03C002C";
end if;
if first_state_sram_input_id = 9699 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 9700 then
	sram_write <= x"03DC0040";
end if;
if first_state_sram_input_id = 9701 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 9702 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 9703 then
	sram_write <= x"82008034";
end if;
if first_state_sram_input_id = 9704 then
	sram_write <= x"07DC0040";
end if;
if first_state_sram_input_id = 9705 then
	sram_write <= x"820097F8";
end if;
if first_state_sram_input_id = 9706 then
	sram_write <= x"C04201DC";
end if;
if first_state_sram_input_id = 9707 then
	sram_write <= x"C8400014";
end if;
if first_state_sram_input_id = 9708 then
	sram_write <= x"C45C0038";
end if;
if first_state_sram_input_id = 9709 then
	sram_write <= x"CC3C0030";
end if;
if first_state_sram_input_id = 9710 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 9711 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 9712 then
	sram_write <= x"03DC0044";
end if;
if first_state_sram_input_id = 9713 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 9714 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 9715 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 9716 then
	sram_write <= x"07DC0044";
end if;
if first_state_sram_input_id = 9717 then
	sram_write <= x"C85C0030";
end if;
if first_state_sram_input_id = 9718 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 9719 then
	sram_write <= x"C03C0038";
end if;
if first_state_sram_input_id = 9720 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 9721 then
	sram_write <= x"03DC0044";
end if;
if first_state_sram_input_id = 9722 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 9723 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 9724 then
	sram_write <= x"82008034";
end if;
if first_state_sram_input_id = 9725 then
	sram_write <= x"07DC0044";
end if;
if first_state_sram_input_id = 9726 then
	sram_write <= x"02800074";
end if;
if first_state_sram_input_id = 9727 then
	sram_write <= x"C03C0028";
end if;
if first_state_sram_input_id = 9728 then
	sram_write <= x"C05C0024";
end if;
if first_state_sram_input_id = 9729 then
	sram_write <= x"C07C0020";
end if;
if first_state_sram_input_id = 9730 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 9731 then
	sram_write <= x"03DC0044";
end if;
if first_state_sram_input_id = 9732 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 9733 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 9734 then
	sram_write <= x"82008280";
end if;
if first_state_sram_input_id = 9735 then
	sram_write <= x"07DC0044";
end if;
if first_state_sram_input_id = 9736 then
	sram_write <= x"C03C0008";
end if;
if first_state_sram_input_id = 9737 then
	sram_write <= x"C0420014";
end if;
if first_state_sram_input_id = 9738 then
	sram_write <= x"C07C0018";
end if;
if first_state_sram_input_id = 9739 then
	sram_write <= x"22860220";
end if;
if first_state_sram_input_id = 9740 then
	sram_write <= x"D0448000";
end if;
if first_state_sram_input_id = 9741 then
	sram_write <= x"C09C001C";
end if;
if first_state_sram_input_id = 9742 then
	sram_write <= x"C8280000";
end if;
if first_state_sram_input_id = 9743 then
	sram_write <= x"CC240000";
end if;
if first_state_sram_input_id = 9744 then
	sram_write <= x"C8280004";
end if;
if first_state_sram_input_id = 9745 then
	sram_write <= x"CC240004";
end if;
if first_state_sram_input_id = 9746 then
	sram_write <= x"C8280008";
end if;
if first_state_sram_input_id = 9747 then
	sram_write <= x"CC240008";
end if;
if first_state_sram_input_id = 9748 then
	sram_write <= x"82009854";
end if;
if first_state_sram_input_id = 9749 then
	sram_write <= x"C05C0018";
end if;
if first_state_sram_input_id = 9750 then
	sram_write <= x"02440001";
end if;
if first_state_sram_input_id = 9751 then
	sram_write <= x"8200952C";
end if;
if first_state_sram_input_id = 9752 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 9753 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 9754 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 9755 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 9756 then
	sram_write <= x"86409C04";
end if;
if first_state_sram_input_id = 9757 then
	sram_write <= x"02800308";
end if;
if first_state_sram_input_id = 9758 then
	sram_write <= x"C8880000";
end if;
if first_state_sram_input_id = 9759 then
	sram_write <= x"02800300";
end if;
if first_state_sram_input_id = 9760 then
	sram_write <= x"C0880000";
end if;
if first_state_sram_input_id = 9761 then
	sram_write <= x"04848000";
end if;
if first_state_sram_input_id = 9762 then
	sram_write <= x"58A80000";
end if;
if first_state_sram_input_id = 9763 then
	sram_write <= x"4888A000";
end if;
if first_state_sram_input_id = 9764 then
	sram_write <= x"02800348";
end if;
if first_state_sram_input_id = 9765 then
	sram_write <= x"02A00324";
end if;
if first_state_sram_input_id = 9766 then
	sram_write <= x"C8AA0000";
end if;
if first_state_sram_input_id = 9767 then
	sram_write <= x"48A8A000";
end if;
if first_state_sram_input_id = 9768 then
	sram_write <= x"40AA2000";
end if;
if first_state_sram_input_id = 9769 then
	sram_write <= x"CCA80000";
end if;
if first_state_sram_input_id = 9770 then
	sram_write <= x"C8AA0004";
end if;
if first_state_sram_input_id = 9771 then
	sram_write <= x"48A8A000";
end if;
if first_state_sram_input_id = 9772 then
	sram_write <= x"40AA4000";
end if;
if first_state_sram_input_id = 9773 then
	sram_write <= x"CCA80004";
end if;
if first_state_sram_input_id = 9774 then
	sram_write <= x"C8AA0008";
end if;
if first_state_sram_input_id = 9775 then
	sram_write <= x"4888A000";
end if;
if first_state_sram_input_id = 9776 then
	sram_write <= x"40886000";
end if;
if first_state_sram_input_id = 9777 then
	sram_write <= x"CC880008";
end if;
if first_state_sram_input_id = 9778 then
	sram_write <= x"02A00000";
end if;
if first_state_sram_input_id = 9779 then
	sram_write <= x"CC7C0000";
end if;
if first_state_sram_input_id = 9780 then
	sram_write <= x"CC5C0008";
end if;
if first_state_sram_input_id = 9781 then
	sram_write <= x"CC3C0010";
end if;
if first_state_sram_input_id = 9782 then
	sram_write <= x"C47C0018";
end if;
if first_state_sram_input_id = 9783 then
	sram_write <= x"C49C001C";
end if;
if first_state_sram_input_id = 9784 then
	sram_write <= x"C43C0020";
end if;
if first_state_sram_input_id = 9785 then
	sram_write <= x"C45C0024";
end if;
if first_state_sram_input_id = 9786 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 9787 then
	sram_write <= x"004A0000";
end if;
if first_state_sram_input_id = 9788 then
	sram_write <= x"00280000";
end if;
if first_state_sram_input_id = 9789 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 9790 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 9791 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 9792 then
	sram_write <= x"8200161C";
end if;
if first_state_sram_input_id = 9793 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 9794 then
	sram_write <= x"022002EC";
end if;
if first_state_sram_input_id = 9795 then
	sram_write <= x"40400000";
end if;
if first_state_sram_input_id = 9796 then
	sram_write <= x"CC020000";
end if;
if first_state_sram_input_id = 9797 then
	sram_write <= x"CC020004";
end if;
if first_state_sram_input_id = 9798 then
	sram_write <= x"CC020008";
end if;
if first_state_sram_input_id = 9799 then
	sram_write <= x"0240030C";
end if;
if first_state_sram_input_id = 9800 then
	sram_write <= x"026001C4";
end if;
if first_state_sram_input_id = 9801 then
	sram_write <= x"C8260000";
end if;
if first_state_sram_input_id = 9802 then
	sram_write <= x"CC240000";
end if;
if first_state_sram_input_id = 9803 then
	sram_write <= x"C8260004";
end if;
if first_state_sram_input_id = 9804 then
	sram_write <= x"CC240004";
end if;
if first_state_sram_input_id = 9805 then
	sram_write <= x"C8260008";
end if;
if first_state_sram_input_id = 9806 then
	sram_write <= x"CC240008";
end if;
if first_state_sram_input_id = 9807 then
	sram_write <= x"02400000";
end if;
if first_state_sram_input_id = 9808 then
	sram_write <= x"C82000A8";
end if;
if first_state_sram_input_id = 9809 then
	sram_write <= x"C07C0024";
end if;
if first_state_sram_input_id = 9810 then
	sram_write <= x"22860220";
end if;
if first_state_sram_input_id = 9811 then
	sram_write <= x"C0BC0020";
end if;
if first_state_sram_input_id = 9812 then
	sram_write <= x"D08A8000";
end if;
if first_state_sram_input_id = 9813 then
	sram_write <= x"C0DC001C";
end if;
if first_state_sram_input_id = 9814 then
	sram_write <= x"C43C0028";
end if;
if first_state_sram_input_id = 9815 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 9816 then
	sram_write <= x"00680000";
end if;
if first_state_sram_input_id = 9817 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 9818 then
	sram_write <= x"004C0000";
end if;
if first_state_sram_input_id = 9819 then
	sram_write <= x"03DC0034";
end if;
if first_state_sram_input_id = 9820 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 9821 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 9822 then
	sram_write <= x"82007A14";
end if;
if first_state_sram_input_id = 9823 then
	sram_write <= x"07DC0034";
end if;
if first_state_sram_input_id = 9824 then
	sram_write <= x"C03C0024";
end if;
if first_state_sram_input_id = 9825 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 9826 then
	sram_write <= x"C07C0020";
end if;
if first_state_sram_input_id = 9827 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 9828 then
	sram_write <= x"C0440000";
end if;
if first_state_sram_input_id = 9829 then
	sram_write <= x"C09C0028";
end if;
if first_state_sram_input_id = 9830 then
	sram_write <= x"C8280000";
end if;
if first_state_sram_input_id = 9831 then
	sram_write <= x"CC240000";
end if;
if first_state_sram_input_id = 9832 then
	sram_write <= x"C8280004";
end if;
if first_state_sram_input_id = 9833 then
	sram_write <= x"CC240004";
end if;
if first_state_sram_input_id = 9834 then
	sram_write <= x"C8280008";
end if;
if first_state_sram_input_id = 9835 then
	sram_write <= x"CC240008";
end if;
if first_state_sram_input_id = 9836 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 9837 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 9838 then
	sram_write <= x"C0440018";
end if;
if first_state_sram_input_id = 9839 then
	sram_write <= x"C09C0018";
end if;
if first_state_sram_input_id = 9840 then
	sram_write <= x"C4840000";
end if;
if first_state_sram_input_id = 9841 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 9842 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 9843 then
	sram_write <= x"C0A40008";
end if;
if first_state_sram_input_id = 9844 then
	sram_write <= x"C0AA0000";
end if;
if first_state_sram_input_id = 9845 then
	sram_write <= x"86A09BCC";
end if;
if first_state_sram_input_id = 9846 then
	sram_write <= x"C0A4000C";
end if;
if first_state_sram_input_id = 9847 then
	sram_write <= x"C0AA0000";
end if;
if first_state_sram_input_id = 9848 then
	sram_write <= x"C45C002C";
end if;
if first_state_sram_input_id = 9849 then
	sram_write <= x"82A09BA8";
end if;
if first_state_sram_input_id = 9850 then
	sram_write <= x"C0A40018";
end if;
if first_state_sram_input_id = 9851 then
	sram_write <= x"C0AA0000";
end if;
if first_state_sram_input_id = 9852 then
	sram_write <= x"02C002E0";
end if;
if first_state_sram_input_id = 9853 then
	sram_write <= x"CC0C0000";
end if;
if first_state_sram_input_id = 9854 then
	sram_write <= x"CC0C0004";
end if;
if first_state_sram_input_id = 9855 then
	sram_write <= x"CC0C0008";
end if;
if first_state_sram_input_id = 9856 then
	sram_write <= x"C0E4001C";
end if;
if first_state_sram_input_id = 9857 then
	sram_write <= x"C1040004";
end if;
if first_state_sram_input_id = 9858 then
	sram_write <= x"03200354";
end if;
if first_state_sram_input_id = 9859 then
	sram_write <= x"22AA0220";
end if;
if first_state_sram_input_id = 9860 then
	sram_write <= x"D0B2A000";
end if;
if first_state_sram_input_id = 9861 then
	sram_write <= x"C0EE0000";
end if;
if first_state_sram_input_id = 9862 then
	sram_write <= x"C1100000";
end if;
if first_state_sram_input_id = 9863 then
	sram_write <= x"03200318";
end if;
if first_state_sram_input_id = 9864 then
	sram_write <= x"C8300000";
end if;
if first_state_sram_input_id = 9865 then
	sram_write <= x"CC320000";
end if;
if first_state_sram_input_id = 9866 then
	sram_write <= x"C8300004";
end if;
if first_state_sram_input_id = 9867 then
	sram_write <= x"CC320004";
end if;
if first_state_sram_input_id = 9868 then
	sram_write <= x"C8300008";
end if;
if first_state_sram_input_id = 9869 then
	sram_write <= x"CC320008";
end if;
if first_state_sram_input_id = 9870 then
	sram_write <= x"032000C4";
end if;
if first_state_sram_input_id = 9871 then
	sram_write <= x"C1320000";
end if;
if first_state_sram_input_id = 9872 then
	sram_write <= x"07320001";
end if;
if first_state_sram_input_id = 9873 then
	sram_write <= x"C4DC0030";
end if;
if first_state_sram_input_id = 9874 then
	sram_write <= x"C51C0034";
end if;
if first_state_sram_input_id = 9875 then
	sram_write <= x"C4FC0038";
end if;
if first_state_sram_input_id = 9876 then
	sram_write <= x"C4BC003C";
end if;
if first_state_sram_input_id = 9877 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 9878 then
	sram_write <= x"00520000";
end if;
if first_state_sram_input_id = 9879 then
	sram_write <= x"00300000";
end if;
if first_state_sram_input_id = 9880 then
	sram_write <= x"03DC0048";
end if;
if first_state_sram_input_id = 9881 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 9882 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 9883 then
	sram_write <= x"8200462C";
end if;
if first_state_sram_input_id = 9884 then
	sram_write <= x"07DC0048";
end if;
if first_state_sram_input_id = 9885 then
	sram_write <= x"C03C003C";
end if;
if first_state_sram_input_id = 9886 then
	sram_write <= x"C04201D8";
end if;
if first_state_sram_input_id = 9887 then
	sram_write <= x"C0640000";
end if;
if first_state_sram_input_id = 9888 then
	sram_write <= x"C8260000";
end if;
if first_state_sram_input_id = 9889 then
	sram_write <= x"C09C0038";
end if;
if first_state_sram_input_id = 9890 then
	sram_write <= x"C8480000";
end if;
if first_state_sram_input_id = 9891 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 9892 then
	sram_write <= x"C8460004";
end if;
if first_state_sram_input_id = 9893 then
	sram_write <= x"C8680004";
end if;
if first_state_sram_input_id = 9894 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 9895 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 9896 then
	sram_write <= x"C8460008";
end if;
if first_state_sram_input_id = 9897 then
	sram_write <= x"C8680008";
end if;
if first_state_sram_input_id = 9898 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 9899 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 9900 then
	sram_write <= x"8E209B04";
end if;
if first_state_sram_input_id = 9901 then
	sram_write <= x"C8400018";
end if;
if first_state_sram_input_id = 9902 then
	sram_write <= x"C45C0040";
end if;
if first_state_sram_input_id = 9903 then
	sram_write <= x"CC3C0048";
end if;
if first_state_sram_input_id = 9904 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 9905 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 9906 then
	sram_write <= x"03DC0058";
end if;
if first_state_sram_input_id = 9907 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 9908 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 9909 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 9910 then
	sram_write <= x"07DC0058";
end if;
if first_state_sram_input_id = 9911 then
	sram_write <= x"C85C0048";
end if;
if first_state_sram_input_id = 9912 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 9913 then
	sram_write <= x"C03C0040";
end if;
if first_state_sram_input_id = 9914 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 9915 then
	sram_write <= x"03DC0058";
end if;
if first_state_sram_input_id = 9916 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 9917 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 9918 then
	sram_write <= x"82008034";
end if;
if first_state_sram_input_id = 9919 then
	sram_write <= x"07DC0058";
end if;
if first_state_sram_input_id = 9920 then
	sram_write <= x"82009B54";
end if;
if first_state_sram_input_id = 9921 then
	sram_write <= x"C04201DC";
end if;
if first_state_sram_input_id = 9922 then
	sram_write <= x"C8400014";
end if;
if first_state_sram_input_id = 9923 then
	sram_write <= x"C45C0050";
end if;
if first_state_sram_input_id = 9924 then
	sram_write <= x"CC3C0048";
end if;
if first_state_sram_input_id = 9925 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 9926 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 9927 then
	sram_write <= x"03DC005C";
end if;
if first_state_sram_input_id = 9928 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 9929 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 9930 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 9931 then
	sram_write <= x"07DC005C";
end if;
if first_state_sram_input_id = 9932 then
	sram_write <= x"C85C0048";
end if;
if first_state_sram_input_id = 9933 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 9934 then
	sram_write <= x"C03C0050";
end if;
if first_state_sram_input_id = 9935 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 9936 then
	sram_write <= x"03DC005C";
end if;
if first_state_sram_input_id = 9937 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 9938 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 9939 then
	sram_write <= x"82008034";
end if;
if first_state_sram_input_id = 9940 then
	sram_write <= x"07DC005C";
end if;
if first_state_sram_input_id = 9941 then
	sram_write <= x"02800074";
end if;
if first_state_sram_input_id = 9942 then
	sram_write <= x"C03C003C";
end if;
if first_state_sram_input_id = 9943 then
	sram_write <= x"C05C0038";
end if;
if first_state_sram_input_id = 9944 then
	sram_write <= x"C07C0034";
end if;
if first_state_sram_input_id = 9945 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 9946 then
	sram_write <= x"03DC005C";
end if;
if first_state_sram_input_id = 9947 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 9948 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 9949 then
	sram_write <= x"82008280";
end if;
if first_state_sram_input_id = 9950 then
	sram_write <= x"07DC005C";
end if;
if first_state_sram_input_id = 9951 then
	sram_write <= x"C03C002C";
end if;
if first_state_sram_input_id = 9952 then
	sram_write <= x"C0420014";
end if;
if first_state_sram_input_id = 9953 then
	sram_write <= x"C0440000";
end if;
if first_state_sram_input_id = 9954 then
	sram_write <= x"C07C0030";
end if;
if first_state_sram_input_id = 9955 then
	sram_write <= x"C8260000";
end if;
if first_state_sram_input_id = 9956 then
	sram_write <= x"CC240000";
end if;
if first_state_sram_input_id = 9957 then
	sram_write <= x"C8260004";
end if;
if first_state_sram_input_id = 9958 then
	sram_write <= x"CC240004";
end if;
if first_state_sram_input_id = 9959 then
	sram_write <= x"C8260008";
end if;
if first_state_sram_input_id = 9960 then
	sram_write <= x"CC240008";
end if;
if first_state_sram_input_id = 9961 then
	sram_write <= x"82009BA8";
end if;
if first_state_sram_input_id = 9962 then
	sram_write <= x"02400001";
end if;
if first_state_sram_input_id = 9963 then
	sram_write <= x"C03C002C";
end if;
if first_state_sram_input_id = 9964 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 9965 then
	sram_write <= x"03DC005C";
end if;
if first_state_sram_input_id = 9966 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 9967 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 9968 then
	sram_write <= x"8200952C";
end if;
if first_state_sram_input_id = 9969 then
	sram_write <= x"07DC005C";
end if;
if first_state_sram_input_id = 9970 then
	sram_write <= x"82009BCC";
end if;
if first_state_sram_input_id = 9971 then
	sram_write <= x"C03C0024";
end if;
if first_state_sram_input_id = 9972 then
	sram_write <= x"06420001";
end if;
if first_state_sram_input_id = 9973 then
	sram_write <= x"C03C0018";
end if;
if first_state_sram_input_id = 9974 then
	sram_write <= x"02220001";
end if;
if first_state_sram_input_id = 9975 then
	sram_write <= x"02600005";
end if;
if first_state_sram_input_id = 9976 then
	sram_write <= x"86269BEC";
end if;
if first_state_sram_input_id = 9977 then
	sram_write <= x"06620005";
end if;
if first_state_sram_input_id = 9978 then
	sram_write <= x"82009BF0";
end if;
if first_state_sram_input_id = 9979 then
	sram_write <= x"00620000";
end if;
if first_state_sram_input_id = 9980 then
	sram_write <= x"C83C0010";
end if;
if first_state_sram_input_id = 9981 then
	sram_write <= x"C85C0008";
end if;
if first_state_sram_input_id = 9982 then
	sram_write <= x"C87C0000";
end if;
if first_state_sram_input_id = 9983 then
	sram_write <= x"C03C0020";
end if;
if first_state_sram_input_id = 9984 then
	sram_write <= x"82009870";
end if;
if first_state_sram_input_id = 9985 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 9986 then
	sram_write <= x"02800308";
end if;
if first_state_sram_input_id = 9987 then
	sram_write <= x"C8280000";
end if;
if first_state_sram_input_id = 9988 then
	sram_write <= x"02800300";
end if;
if first_state_sram_input_id = 9989 then
	sram_write <= x"C0880004";
end if;
if first_state_sram_input_id = 9990 then
	sram_write <= x"04448000";
end if;
if first_state_sram_input_id = 9991 then
	sram_write <= x"58440000";
end if;
if first_state_sram_input_id = 9992 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 9993 then
	sram_write <= x"02400330";
end if;
if first_state_sram_input_id = 9994 then
	sram_write <= x"C8440000";
end if;
if first_state_sram_input_id = 9995 then
	sram_write <= x"48424000";
end if;
if first_state_sram_input_id = 9996 then
	sram_write <= x"0280033C";
end if;
if first_state_sram_input_id = 9997 then
	sram_write <= x"C8680000";
end if;
if first_state_sram_input_id = 9998 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 9999 then
	sram_write <= x"C8640004";
end if;
if first_state_sram_input_id = 10000 then
	sram_write <= x"48626000";
end if;
if first_state_sram_input_id = 10001 then
	sram_write <= x"C8880004";
end if;
if first_state_sram_input_id = 10002 then
	sram_write <= x"40668000";
end if;
if first_state_sram_input_id = 10003 then
	sram_write <= x"C8840008";
end if;
if first_state_sram_input_id = 10004 then
	sram_write <= x"48228000";
end if;
if first_state_sram_input_id = 10005 then
	sram_write <= x"C8880008";
end if;
if first_state_sram_input_id = 10006 then
	sram_write <= x"40228000";
end if;
if first_state_sram_input_id = 10007 then
	sram_write <= x"024002F8";
end if;
if first_state_sram_input_id = 10008 then
	sram_write <= x"C0440000";
end if;
if first_state_sram_input_id = 10009 then
	sram_write <= x"06440001";
end if;
if first_state_sram_input_id = 10010 then
	sram_write <= x"41E06000";
end if;
if first_state_sram_input_id = 10011 then
	sram_write <= x"40602000";
end if;
if first_state_sram_input_id = 10012 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 10013 then
	sram_write <= x"4041E000";
end if;
if first_state_sram_input_id = 10014 then
	sram_write <= x"82009870";
end if;
if first_state_sram_input_id = 10015 then
	sram_write <= x"02C002F8";
end if;
if first_state_sram_input_id = 10016 then
	sram_write <= x"C0EC0000";
end if;
if first_state_sram_input_id = 10017 then
	sram_write <= x"862E9C8C";
end if;
if first_state_sram_input_id = 10018 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 10019 then
	sram_write <= x"02E002EC";
end if;
if first_state_sram_input_id = 10020 then
	sram_write <= x"23020220";
end if;
if first_state_sram_input_id = 10021 then
	sram_write <= x"D1090000";
end if;
if first_state_sram_input_id = 10022 then
	sram_write <= x"C1100000";
end if;
if first_state_sram_input_id = 10023 then
	sram_write <= x"C8300000";
end if;
if first_state_sram_input_id = 10024 then
	sram_write <= x"CC2E0000";
end if;
if first_state_sram_input_id = 10025 then
	sram_write <= x"C8300004";
end if;
if first_state_sram_input_id = 10026 then
	sram_write <= x"CC2E0004";
end if;
if first_state_sram_input_id = 10027 then
	sram_write <= x"C8300008";
end if;
if first_state_sram_input_id = 10028 then
	sram_write <= x"CC2E0008";
end if;
if first_state_sram_input_id = 10029 then
	sram_write <= x"03040001";
end if;
if first_state_sram_input_id = 10030 then
	sram_write <= x"C12C0004";
end if;
if first_state_sram_input_id = 10031 then
	sram_write <= x"87129CC8";
end if;
if first_state_sram_input_id = 10032 then
	sram_write <= x"03000000";
end if;
if first_state_sram_input_id = 10033 then
	sram_write <= x"82009CF8";
end if;
if first_state_sram_input_id = 10034 then
	sram_write <= x"86049CD4";
end if;
if first_state_sram_input_id = 10035 then
	sram_write <= x"03000000";
end if;
if first_state_sram_input_id = 10036 then
	sram_write <= x"82009CF8";
end if;
if first_state_sram_input_id = 10037 then
	sram_write <= x"03020001";
end if;
if first_state_sram_input_id = 10038 then
	sram_write <= x"C12C0000";
end if;
if first_state_sram_input_id = 10039 then
	sram_write <= x"87129CE8";
end if;
if first_state_sram_input_id = 10040 then
	sram_write <= x"03000000";
end if;
if first_state_sram_input_id = 10041 then
	sram_write <= x"82009CF8";
end if;
if first_state_sram_input_id = 10042 then
	sram_write <= x"86029CF4";
end if;
if first_state_sram_input_id = 10043 then
	sram_write <= x"03000000";
end if;
if first_state_sram_input_id = 10044 then
	sram_write <= x"82009CF8";
end if;
if first_state_sram_input_id = 10045 then
	sram_write <= x"03000001";
end if;
if first_state_sram_input_id = 10046 then
	sram_write <= x"C4BC0000";
end if;
if first_state_sram_input_id = 10047 then
	sram_write <= x"C47C0004";
end if;
if first_state_sram_input_id = 10048 then
	sram_write <= x"C45C0008";
end if;
if first_state_sram_input_id = 10049 then
	sram_write <= x"C49C000C";
end if;
if first_state_sram_input_id = 10050 then
	sram_write <= x"C4DC0010";
end if;
if first_state_sram_input_id = 10051 then
	sram_write <= x"C43C0014";
end if;
if first_state_sram_input_id = 10052 then
	sram_write <= x"C4FC0018";
end if;
if first_state_sram_input_id = 10053 then
	sram_write <= x"83009E4C";
end if;
if first_state_sram_input_id = 10054 then
	sram_write <= x"03000000";
end if;
if first_state_sram_input_id = 10055 then
	sram_write <= x"23220220";
end if;
if first_state_sram_input_id = 10056 then
	sram_write <= x"D1292000";
end if;
if first_state_sram_input_id = 10057 then
	sram_write <= x"C1520008";
end if;
if first_state_sram_input_id = 10058 then
	sram_write <= x"C1540000";
end if;
if first_state_sram_input_id = 10059 then
	sram_write <= x"87409E48";
end if;
if first_state_sram_input_id = 10060 then
	sram_write <= x"C1520008";
end if;
if first_state_sram_input_id = 10061 then
	sram_write <= x"C1540000";
end if;
if first_state_sram_input_id = 10062 then
	sram_write <= x"22C20220";
end if;
if first_state_sram_input_id = 10063 then
	sram_write <= x"D0C6C000";
end if;
if first_state_sram_input_id = 10064 then
	sram_write <= x"C0CC0008";
end if;
if first_state_sram_input_id = 10065 then
	sram_write <= x"C0CC0000";
end if;
if first_state_sram_input_id = 10066 then
	sram_write <= x"82D49D54";
end if;
if first_state_sram_input_id = 10067 then
	sram_write <= x"02C00000";
end if;
if first_state_sram_input_id = 10068 then
	sram_write <= x"82009DB4";
end if;
if first_state_sram_input_id = 10069 then
	sram_write <= x"22C20220";
end if;
if first_state_sram_input_id = 10070 then
	sram_write <= x"D0CAC000";
end if;
if first_state_sram_input_id = 10071 then
	sram_write <= x"C0CC0008";
end if;
if first_state_sram_input_id = 10072 then
	sram_write <= x"C0CC0000";
end if;
if first_state_sram_input_id = 10073 then
	sram_write <= x"82D49D70";
end if;
if first_state_sram_input_id = 10074 then
	sram_write <= x"02C00000";
end if;
if first_state_sram_input_id = 10075 then
	sram_write <= x"82009DB4";
end if;
if first_state_sram_input_id = 10076 then
	sram_write <= x"06C20001";
end if;
if first_state_sram_input_id = 10077 then
	sram_write <= x"22CC0220";
end if;
if first_state_sram_input_id = 10078 then
	sram_write <= x"D0C8C000";
end if;
if first_state_sram_input_id = 10079 then
	sram_write <= x"C0CC0008";
end if;
if first_state_sram_input_id = 10080 then
	sram_write <= x"C0CC0000";
end if;
if first_state_sram_input_id = 10081 then
	sram_write <= x"82D49D90";
end if;
if first_state_sram_input_id = 10082 then
	sram_write <= x"02C00000";
end if;
if first_state_sram_input_id = 10083 then
	sram_write <= x"82009DB4";
end if;
if first_state_sram_input_id = 10084 then
	sram_write <= x"02C20001";
end if;
if first_state_sram_input_id = 10085 then
	sram_write <= x"22CC0220";
end if;
if first_state_sram_input_id = 10086 then
	sram_write <= x"D0C8C000";
end if;
if first_state_sram_input_id = 10087 then
	sram_write <= x"C0CC0008";
end if;
if first_state_sram_input_id = 10088 then
	sram_write <= x"C0CC0000";
end if;
if first_state_sram_input_id = 10089 then
	sram_write <= x"82D49DB0";
end if;
if first_state_sram_input_id = 10090 then
	sram_write <= x"02C00000";
end if;
if first_state_sram_input_id = 10091 then
	sram_write <= x"82009DB4";
end if;
if first_state_sram_input_id = 10092 then
	sram_write <= x"02C00001";
end if;
if first_state_sram_input_id = 10093 then
	sram_write <= x"82C09E24";
end if;
if first_state_sram_input_id = 10094 then
	sram_write <= x"C0D2000C";
end if;
if first_state_sram_input_id = 10095 then
	sram_write <= x"C0CC0000";
end if;
if first_state_sram_input_id = 10096 then
	sram_write <= x"82C09DF0";
end if;
if first_state_sram_input_id = 10097 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10098 then
	sram_write <= x"00460000";
end if;
if first_state_sram_input_id = 10099 then
	sram_write <= x"00680000";
end if;
if first_state_sram_input_id = 10100 then
	sram_write <= x"008A0000";
end if;
if first_state_sram_input_id = 10101 then
	sram_write <= x"00B00000";
end if;
if first_state_sram_input_id = 10102 then
	sram_write <= x"03DC0024";
end if;
if first_state_sram_input_id = 10103 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10104 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10105 then
	sram_write <= x"82008F34";
end if;
if first_state_sram_input_id = 10106 then
	sram_write <= x"07DC0024";
end if;
if first_state_sram_input_id = 10107 then
	sram_write <= x"82009DF0";
end if;
if first_state_sram_input_id = 10108 then
	sram_write <= x"02C00001";
end if;
if first_state_sram_input_id = 10109 then
	sram_write <= x"C03C0014";
end if;
if first_state_sram_input_id = 10110 then
	sram_write <= x"C05C0008";
end if;
if first_state_sram_input_id = 10111 then
	sram_write <= x"C07C0004";
end if;
if first_state_sram_input_id = 10112 then
	sram_write <= x"C09C000C";
end if;
if first_state_sram_input_id = 10113 then
	sram_write <= x"C0BC0000";
end if;
if first_state_sram_input_id = 10114 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10115 then
	sram_write <= x"03DC0024";
end if;
if first_state_sram_input_id = 10116 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10117 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10118 then
	sram_write <= x"8200925C";
end if;
if first_state_sram_input_id = 10119 then
	sram_write <= x"07DC0024";
end if;
if first_state_sram_input_id = 10120 then
	sram_write <= x"82009E44";
end if;
if first_state_sram_input_id = 10121 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10122 then
	sram_write <= x"00500000";
end if;
if first_state_sram_input_id = 10123 then
	sram_write <= x"00320000";
end if;
if first_state_sram_input_id = 10124 then
	sram_write <= x"03DC0024";
end if;
if first_state_sram_input_id = 10125 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10126 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10127 then
	sram_write <= x"820090E0";
end if;
if first_state_sram_input_id = 10128 then
	sram_write <= x"07DC0024";
end if;
if first_state_sram_input_id = 10129 then
	sram_write <= x"82009E48";
end if;
if first_state_sram_input_id = 10130 then
	sram_write <= x"82009EBC";
end if;
if first_state_sram_input_id = 10131 then
	sram_write <= x"23020220";
end if;
if first_state_sram_input_id = 10132 then
	sram_write <= x"D1090000";
end if;
if first_state_sram_input_id = 10133 then
	sram_write <= x"03200000";
end if;
if first_state_sram_input_id = 10134 then
	sram_write <= x"C1500008";
end if;
if first_state_sram_input_id = 10135 then
	sram_write <= x"C1540000";
end if;
if first_state_sram_input_id = 10136 then
	sram_write <= x"87409EBC";
end if;
if first_state_sram_input_id = 10137 then
	sram_write <= x"C150000C";
end if;
if first_state_sram_input_id = 10138 then
	sram_write <= x"C1540000";
end if;
if first_state_sram_input_id = 10139 then
	sram_write <= x"C51C001C";
end if;
if first_state_sram_input_id = 10140 then
	sram_write <= x"83409E98";
end if;
if first_state_sram_input_id = 10141 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10142 then
	sram_write <= x"00520000";
end if;
if first_state_sram_input_id = 10143 then
	sram_write <= x"00300000";
end if;
if first_state_sram_input_id = 10144 then
	sram_write <= x"03DC0028";
end if;
if first_state_sram_input_id = 10145 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10146 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10147 then
	sram_write <= x"8200874C";
end if;
if first_state_sram_input_id = 10148 then
	sram_write <= x"07DC0028";
end if;
if first_state_sram_input_id = 10149 then
	sram_write <= x"82009E98";
end if;
if first_state_sram_input_id = 10150 then
	sram_write <= x"02400001";
end if;
if first_state_sram_input_id = 10151 then
	sram_write <= x"C03C001C";
end if;
if first_state_sram_input_id = 10152 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10153 then
	sram_write <= x"03DC0028";
end if;
if first_state_sram_input_id = 10154 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10155 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10156 then
	sram_write <= x"820090E0";
end if;
if first_state_sram_input_id = 10157 then
	sram_write <= x"07DC0028";
end if;
if first_state_sram_input_id = 10158 then
	sram_write <= x"82009EBC";
end if;
if first_state_sram_input_id = 10159 then
	sram_write <= x"C03C0018";
end if;
if first_state_sram_input_id = 10160 then
	sram_write <= x"C8220000";
end if;
if first_state_sram_input_id = 10161 then
	sram_write <= x"54420000";
end if;
if first_state_sram_input_id = 10162 then
	sram_write <= x"026000FF";
end if;
if first_state_sram_input_id = 10163 then
	sram_write <= x"86649EE0";
end if;
if first_state_sram_input_id = 10164 then
	sram_write <= x"86409ED8";
end if;
if first_state_sram_input_id = 10165 then
	sram_write <= x"82009EDC";
end if;
if first_state_sram_input_id = 10166 then
	sram_write <= x"02400000";
end if;
if first_state_sram_input_id = 10167 then
	sram_write <= x"82009EE4";
end if;
if first_state_sram_input_id = 10168 then
	sram_write <= x"024000FF";
end if;
if first_state_sram_input_id = 10169 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10170 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 10171 then
	sram_write <= x"03DC0028";
end if;
if first_state_sram_input_id = 10172 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10173 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10174 then
	sram_write <= x"8200078C";
end if;
if first_state_sram_input_id = 10175 then
	sram_write <= x"07DC0028";
end if;
if first_state_sram_input_id = 10176 then
	sram_write <= x"C03C0018";
end if;
if first_state_sram_input_id = 10177 then
	sram_write <= x"C8220004";
end if;
if first_state_sram_input_id = 10178 then
	sram_write <= x"54420000";
end if;
if first_state_sram_input_id = 10179 then
	sram_write <= x"026000FF";
end if;
if first_state_sram_input_id = 10180 then
	sram_write <= x"86649F24";
end if;
if first_state_sram_input_id = 10181 then
	sram_write <= x"86409F1C";
end if;
if first_state_sram_input_id = 10182 then
	sram_write <= x"82009F20";
end if;
if first_state_sram_input_id = 10183 then
	sram_write <= x"02400000";
end if;
if first_state_sram_input_id = 10184 then
	sram_write <= x"82009F28";
end if;
if first_state_sram_input_id = 10185 then
	sram_write <= x"024000FF";
end if;
if first_state_sram_input_id = 10186 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10187 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 10188 then
	sram_write <= x"03DC0028";
end if;
if first_state_sram_input_id = 10189 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10190 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10191 then
	sram_write <= x"8200078C";
end if;
if first_state_sram_input_id = 10192 then
	sram_write <= x"07DC0028";
end if;
if first_state_sram_input_id = 10193 then
	sram_write <= x"C03C0018";
end if;
if first_state_sram_input_id = 10194 then
	sram_write <= x"C8220008";
end if;
if first_state_sram_input_id = 10195 then
	sram_write <= x"54420000";
end if;
if first_state_sram_input_id = 10196 then
	sram_write <= x"026000FF";
end if;
if first_state_sram_input_id = 10197 then
	sram_write <= x"86649F68";
end if;
if first_state_sram_input_id = 10198 then
	sram_write <= x"86409F60";
end if;
if first_state_sram_input_id = 10199 then
	sram_write <= x"82009F64";
end if;
if first_state_sram_input_id = 10200 then
	sram_write <= x"02400000";
end if;
if first_state_sram_input_id = 10201 then
	sram_write <= x"82009F6C";
end if;
if first_state_sram_input_id = 10202 then
	sram_write <= x"024000FF";
end if;
if first_state_sram_input_id = 10203 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10204 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 10205 then
	sram_write <= x"03DC0028";
end if;
if first_state_sram_input_id = 10206 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10207 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10208 then
	sram_write <= x"8200078C";
end if;
if first_state_sram_input_id = 10209 then
	sram_write <= x"07DC0028";
end if;
if first_state_sram_input_id = 10210 then
	sram_write <= x"C03C0014";
end if;
if first_state_sram_input_id = 10211 then
	sram_write <= x"02220001";
end if;
if first_state_sram_input_id = 10212 then
	sram_write <= x"C05C0010";
end if;
if first_state_sram_input_id = 10213 then
	sram_write <= x"C0640000";
end if;
if first_state_sram_input_id = 10214 then
	sram_write <= x"86269FA0";
end if;
if first_state_sram_input_id = 10215 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 10216 then
	sram_write <= x"22620220";
end if;
if first_state_sram_input_id = 10217 then
	sram_write <= x"C09C000C";
end if;
if first_state_sram_input_id = 10218 then
	sram_write <= x"D0686000";
end if;
if first_state_sram_input_id = 10219 then
	sram_write <= x"C0660000";
end if;
if first_state_sram_input_id = 10220 then
	sram_write <= x"C8260000";
end if;
if first_state_sram_input_id = 10221 then
	sram_write <= x"C0BC0018";
end if;
if first_state_sram_input_id = 10222 then
	sram_write <= x"CC2A0000";
end if;
if first_state_sram_input_id = 10223 then
	sram_write <= x"C8260004";
end if;
if first_state_sram_input_id = 10224 then
	sram_write <= x"CC2A0004";
end if;
if first_state_sram_input_id = 10225 then
	sram_write <= x"C8260008";
end if;
if first_state_sram_input_id = 10226 then
	sram_write <= x"CC2A0008";
end if;
if first_state_sram_input_id = 10227 then
	sram_write <= x"C07C0008";
end if;
if first_state_sram_input_id = 10228 then
	sram_write <= x"02C60001";
end if;
if first_state_sram_input_id = 10229 then
	sram_write <= x"C0E40004";
end if;
if first_state_sram_input_id = 10230 then
	sram_write <= x"86CE9FE4";
end if;
if first_state_sram_input_id = 10231 then
	sram_write <= x"02400000";
end if;
if first_state_sram_input_id = 10232 then
	sram_write <= x"8200A014";
end if;
if first_state_sram_input_id = 10233 then
	sram_write <= x"86069FF0";
end if;
if first_state_sram_input_id = 10234 then
	sram_write <= x"02400000";
end if;
if first_state_sram_input_id = 10235 then
	sram_write <= x"8200A014";
end if;
if first_state_sram_input_id = 10236 then
	sram_write <= x"02C20001";
end if;
if first_state_sram_input_id = 10237 then
	sram_write <= x"C0440000";
end if;
if first_state_sram_input_id = 10238 then
	sram_write <= x"86C4A004";
end if;
if first_state_sram_input_id = 10239 then
	sram_write <= x"02400000";
end if;
if first_state_sram_input_id = 10240 then
	sram_write <= x"8200A014";
end if;
if first_state_sram_input_id = 10241 then
	sram_write <= x"8602A010";
end if;
if first_state_sram_input_id = 10242 then
	sram_write <= x"02400000";
end if;
if first_state_sram_input_id = 10243 then
	sram_write <= x"8200A014";
end if;
if first_state_sram_input_id = 10244 then
	sram_write <= x"02400001";
end if;
if first_state_sram_input_id = 10245 then
	sram_write <= x"C43C0020";
end if;
if first_state_sram_input_id = 10246 then
	sram_write <= x"8240A054";
end if;
if first_state_sram_input_id = 10247 then
	sram_write <= x"02C00000";
end if;
if first_state_sram_input_id = 10248 then
	sram_write <= x"C05C0004";
end if;
if first_state_sram_input_id = 10249 then
	sram_write <= x"C0FC0000";
end if;
if first_state_sram_input_id = 10250 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10251 then
	sram_write <= x"00AE0000";
end if;
if first_state_sram_input_id = 10252 then
	sram_write <= x"01260000";
end if;
if first_state_sram_input_id = 10253 then
	sram_write <= x"00640000";
end if;
if first_state_sram_input_id = 10254 then
	sram_write <= x"00520000";
end if;
if first_state_sram_input_id = 10255 then
	sram_write <= x"03DC002C";
end if;
if first_state_sram_input_id = 10256 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10257 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10258 then
	sram_write <= x"8200925C";
end if;
if first_state_sram_input_id = 10259 then
	sram_write <= x"07DC002C";
end if;
if first_state_sram_input_id = 10260 then
	sram_write <= x"8200A080";
end if;
if first_state_sram_input_id = 10261 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 10262 then
	sram_write <= x"D0484000";
end if;
if first_state_sram_input_id = 10263 then
	sram_write <= x"02C00000";
end if;
if first_state_sram_input_id = 10264 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10265 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 10266 then
	sram_write <= x"004C0000";
end if;
if first_state_sram_input_id = 10267 then
	sram_write <= x"03DC002C";
end if;
if first_state_sram_input_id = 10268 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10269 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10270 then
	sram_write <= x"820090E0";
end if;
if first_state_sram_input_id = 10271 then
	sram_write <= x"07DC002C";
end if;
if first_state_sram_input_id = 10272 then
	sram_write <= x"C03C0018";
end if;
if first_state_sram_input_id = 10273 then
	sram_write <= x"C8220000";
end if;
if first_state_sram_input_id = 10274 then
	sram_write <= x"54420000";
end if;
if first_state_sram_input_id = 10275 then
	sram_write <= x"026000FF";
end if;
if first_state_sram_input_id = 10276 then
	sram_write <= x"8664A0A4";
end if;
if first_state_sram_input_id = 10277 then
	sram_write <= x"8640A09C";
end if;
if first_state_sram_input_id = 10278 then
	sram_write <= x"8200A0A0";
end if;
if first_state_sram_input_id = 10279 then
	sram_write <= x"02400000";
end if;
if first_state_sram_input_id = 10280 then
	sram_write <= x"8200A0A8";
end if;
if first_state_sram_input_id = 10281 then
	sram_write <= x"024000FF";
end if;
if first_state_sram_input_id = 10282 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10283 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 10284 then
	sram_write <= x"03DC002C";
end if;
if first_state_sram_input_id = 10285 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10286 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10287 then
	sram_write <= x"8200078C";
end if;
if first_state_sram_input_id = 10288 then
	sram_write <= x"07DC002C";
end if;
if first_state_sram_input_id = 10289 then
	sram_write <= x"C03C0018";
end if;
if first_state_sram_input_id = 10290 then
	sram_write <= x"C8220004";
end if;
if first_state_sram_input_id = 10291 then
	sram_write <= x"54420000";
end if;
if first_state_sram_input_id = 10292 then
	sram_write <= x"026000FF";
end if;
if first_state_sram_input_id = 10293 then
	sram_write <= x"8664A0E8";
end if;
if first_state_sram_input_id = 10294 then
	sram_write <= x"8640A0E0";
end if;
if first_state_sram_input_id = 10295 then
	sram_write <= x"8200A0E4";
end if;
if first_state_sram_input_id = 10296 then
	sram_write <= x"02400000";
end if;
if first_state_sram_input_id = 10297 then
	sram_write <= x"8200A0EC";
end if;
if first_state_sram_input_id = 10298 then
	sram_write <= x"024000FF";
end if;
if first_state_sram_input_id = 10299 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10300 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 10301 then
	sram_write <= x"03DC002C";
end if;
if first_state_sram_input_id = 10302 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10303 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10304 then
	sram_write <= x"8200078C";
end if;
if first_state_sram_input_id = 10305 then
	sram_write <= x"07DC002C";
end if;
if first_state_sram_input_id = 10306 then
	sram_write <= x"C03C0018";
end if;
if first_state_sram_input_id = 10307 then
	sram_write <= x"C8220008";
end if;
if first_state_sram_input_id = 10308 then
	sram_write <= x"54220000";
end if;
if first_state_sram_input_id = 10309 then
	sram_write <= x"024000FF";
end if;
if first_state_sram_input_id = 10310 then
	sram_write <= x"8642A12C";
end if;
if first_state_sram_input_id = 10311 then
	sram_write <= x"8620A124";
end if;
if first_state_sram_input_id = 10312 then
	sram_write <= x"8200A128";
end if;
if first_state_sram_input_id = 10313 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 10314 then
	sram_write <= x"8200A130";
end if;
if first_state_sram_input_id = 10315 then
	sram_write <= x"022000FF";
end if;
if first_state_sram_input_id = 10316 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10317 then
	sram_write <= x"03DC002C";
end if;
if first_state_sram_input_id = 10318 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10319 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10320 then
	sram_write <= x"8200078C";
end if;
if first_state_sram_input_id = 10321 then
	sram_write <= x"07DC002C";
end if;
if first_state_sram_input_id = 10322 then
	sram_write <= x"C03C0020";
end if;
if first_state_sram_input_id = 10323 then
	sram_write <= x"02220001";
end if;
if first_state_sram_input_id = 10324 then
	sram_write <= x"C05C0008";
end if;
if first_state_sram_input_id = 10325 then
	sram_write <= x"C07C0004";
end if;
if first_state_sram_input_id = 10326 then
	sram_write <= x"C09C000C";
end if;
if first_state_sram_input_id = 10327 then
	sram_write <= x"C0BC0000";
end if;
if first_state_sram_input_id = 10328 then
	sram_write <= x"82009C7C";
end if;
if first_state_sram_input_id = 10329 then
	sram_write <= x"02C002F8";
end if;
if first_state_sram_input_id = 10330 then
	sram_write <= x"C0EC0004";
end if;
if first_state_sram_input_id = 10331 then
	sram_write <= x"862EA174";
end if;
if first_state_sram_input_id = 10332 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 10333 then
	sram_write <= x"C0EC0004";
end if;
if first_state_sram_input_id = 10334 then
	sram_write <= x"06EE0001";
end if;
if first_state_sram_input_id = 10335 then
	sram_write <= x"C4BC0000";
end if;
if first_state_sram_input_id = 10336 then
	sram_write <= x"C49C0004";
end if;
if first_state_sram_input_id = 10337 then
	sram_write <= x"C45C0008";
end if;
if first_state_sram_input_id = 10338 then
	sram_write <= x"C43C000C";
end if;
if first_state_sram_input_id = 10339 then
	sram_write <= x"C47C0010";
end if;
if first_state_sram_input_id = 10340 then
	sram_write <= x"C4DC0014";
end if;
if first_state_sram_input_id = 10341 then
	sram_write <= x"862EA19C";
end if;
if first_state_sram_input_id = 10342 then
	sram_write <= x"8200A1C4";
end if;
if first_state_sram_input_id = 10343 then
	sram_write <= x"02E20001";
end if;
if first_state_sram_input_id = 10344 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10345 then
	sram_write <= x"006A0000";
end if;
if first_state_sram_input_id = 10346 then
	sram_write <= x"004E0000";
end if;
if first_state_sram_input_id = 10347 then
	sram_write <= x"00280000";
end if;
if first_state_sram_input_id = 10348 then
	sram_write <= x"03DC0020";
end if;
if first_state_sram_input_id = 10349 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10350 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10351 then
	sram_write <= x"82009C08";
end if;
if first_state_sram_input_id = 10352 then
	sram_write <= x"07DC0020";
end if;
if first_state_sram_input_id = 10353 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 10354 then
	sram_write <= x"C05C0014";
end if;
if first_state_sram_input_id = 10355 then
	sram_write <= x"C0640000";
end if;
if first_state_sram_input_id = 10356 then
	sram_write <= x"8606A1D8";
end if;
if first_state_sram_input_id = 10357 then
	sram_write <= x"8200A390";
end if;
if first_state_sram_input_id = 10358 then
	sram_write <= x"026002EC";
end if;
if first_state_sram_input_id = 10359 then
	sram_write <= x"C09C0010";
end if;
if first_state_sram_input_id = 10360 then
	sram_write <= x"C0A80000";
end if;
if first_state_sram_input_id = 10361 then
	sram_write <= x"C0AA0000";
end if;
if first_state_sram_input_id = 10362 then
	sram_write <= x"C82A0000";
end if;
if first_state_sram_input_id = 10363 then
	sram_write <= x"CC260000";
end if;
if first_state_sram_input_id = 10364 then
	sram_write <= x"C82A0004";
end if;
if first_state_sram_input_id = 10365 then
	sram_write <= x"CC260004";
end if;
if first_state_sram_input_id = 10366 then
	sram_write <= x"C82A0008";
end if;
if first_state_sram_input_id = 10367 then
	sram_write <= x"CC260008";
end if;
if first_state_sram_input_id = 10368 then
	sram_write <= x"C0BC000C";
end if;
if first_state_sram_input_id = 10369 then
	sram_write <= x"02CA0001";
end if;
if first_state_sram_input_id = 10370 then
	sram_write <= x"C0E40004";
end if;
if first_state_sram_input_id = 10371 then
	sram_write <= x"86CEA218";
end if;
if first_state_sram_input_id = 10372 then
	sram_write <= x"02C00000";
end if;
if first_state_sram_input_id = 10373 then
	sram_write <= x"8200A23C";
end if;
if first_state_sram_input_id = 10374 then
	sram_write <= x"860AA224";
end if;
if first_state_sram_input_id = 10375 then
	sram_write <= x"02C00000";
end if;
if first_state_sram_input_id = 10376 then
	sram_write <= x"8200A23C";
end if;
if first_state_sram_input_id = 10377 then
	sram_write <= x"02C00001";
end if;
if first_state_sram_input_id = 10378 then
	sram_write <= x"C0E40000";
end if;
if first_state_sram_input_id = 10379 then
	sram_write <= x"86CEA238";
end if;
if first_state_sram_input_id = 10380 then
	sram_write <= x"02C00000";
end if;
if first_state_sram_input_id = 10381 then
	sram_write <= x"8200A23C";
end if;
if first_state_sram_input_id = 10382 then
	sram_write <= x"02C00001";
end if;
if first_state_sram_input_id = 10383 then
	sram_write <= x"C47C0018";
end if;
if first_state_sram_input_id = 10384 then
	sram_write <= x"82C0A278";
end if;
if first_state_sram_input_id = 10385 then
	sram_write <= x"02C00000";
end if;
if first_state_sram_input_id = 10386 then
	sram_write <= x"C0FC0008";
end if;
if first_state_sram_input_id = 10387 then
	sram_write <= x"C11C0004";
end if;
if first_state_sram_input_id = 10388 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10389 then
	sram_write <= x"006E0000";
end if;
if first_state_sram_input_id = 10390 then
	sram_write <= x"004A0000";
end if;
if first_state_sram_input_id = 10391 then
	sram_write <= x"00B00000";
end if;
if first_state_sram_input_id = 10392 then
	sram_write <= x"03DC0024";
end if;
if first_state_sram_input_id = 10393 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10394 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10395 then
	sram_write <= x"8200925C";
end if;
if first_state_sram_input_id = 10396 then
	sram_write <= x"07DC0024";
end if;
if first_state_sram_input_id = 10397 then
	sram_write <= x"8200A29C";
end if;
if first_state_sram_input_id = 10398 then
	sram_write <= x"C0280000";
end if;
if first_state_sram_input_id = 10399 then
	sram_write <= x"02C00000";
end if;
if first_state_sram_input_id = 10400 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10401 then
	sram_write <= x"004C0000";
end if;
if first_state_sram_input_id = 10402 then
	sram_write <= x"03DC0024";
end if;
if first_state_sram_input_id = 10403 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10404 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10405 then
	sram_write <= x"820090E0";
end if;
if first_state_sram_input_id = 10406 then
	sram_write <= x"07DC0024";
end if;
if first_state_sram_input_id = 10407 then
	sram_write <= x"C03C0018";
end if;
if first_state_sram_input_id = 10408 then
	sram_write <= x"C8220000";
end if;
if first_state_sram_input_id = 10409 then
	sram_write <= x"54420000";
end if;
if first_state_sram_input_id = 10410 then
	sram_write <= x"026000FF";
end if;
if first_state_sram_input_id = 10411 then
	sram_write <= x"8664A2C0";
end if;
if first_state_sram_input_id = 10412 then
	sram_write <= x"8640A2B8";
end if;
if first_state_sram_input_id = 10413 then
	sram_write <= x"8200A2BC";
end if;
if first_state_sram_input_id = 10414 then
	sram_write <= x"02400000";
end if;
if first_state_sram_input_id = 10415 then
	sram_write <= x"8200A2C4";
end if;
if first_state_sram_input_id = 10416 then
	sram_write <= x"024000FF";
end if;
if first_state_sram_input_id = 10417 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10418 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 10419 then
	sram_write <= x"03DC0024";
end if;
if first_state_sram_input_id = 10420 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10421 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10422 then
	sram_write <= x"8200078C";
end if;
if first_state_sram_input_id = 10423 then
	sram_write <= x"07DC0024";
end if;
if first_state_sram_input_id = 10424 then
	sram_write <= x"C03C0018";
end if;
if first_state_sram_input_id = 10425 then
	sram_write <= x"C8220004";
end if;
if first_state_sram_input_id = 10426 then
	sram_write <= x"54420000";
end if;
if first_state_sram_input_id = 10427 then
	sram_write <= x"026000FF";
end if;
if first_state_sram_input_id = 10428 then
	sram_write <= x"8664A304";
end if;
if first_state_sram_input_id = 10429 then
	sram_write <= x"8640A2FC";
end if;
if first_state_sram_input_id = 10430 then
	sram_write <= x"8200A300";
end if;
if first_state_sram_input_id = 10431 then
	sram_write <= x"02400000";
end if;
if first_state_sram_input_id = 10432 then
	sram_write <= x"8200A308";
end if;
if first_state_sram_input_id = 10433 then
	sram_write <= x"024000FF";
end if;
if first_state_sram_input_id = 10434 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10435 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 10436 then
	sram_write <= x"03DC0024";
end if;
if first_state_sram_input_id = 10437 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10438 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10439 then
	sram_write <= x"8200078C";
end if;
if first_state_sram_input_id = 10440 then
	sram_write <= x"07DC0024";
end if;
if first_state_sram_input_id = 10441 then
	sram_write <= x"C03C0018";
end if;
if first_state_sram_input_id = 10442 then
	sram_write <= x"C8220008";
end if;
if first_state_sram_input_id = 10443 then
	sram_write <= x"54220000";
end if;
if first_state_sram_input_id = 10444 then
	sram_write <= x"024000FF";
end if;
if first_state_sram_input_id = 10445 then
	sram_write <= x"8642A348";
end if;
if first_state_sram_input_id = 10446 then
	sram_write <= x"8620A340";
end if;
if first_state_sram_input_id = 10447 then
	sram_write <= x"8200A344";
end if;
if first_state_sram_input_id = 10448 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 10449 then
	sram_write <= x"8200A34C";
end if;
if first_state_sram_input_id = 10450 then
	sram_write <= x"022000FF";
end if;
if first_state_sram_input_id = 10451 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10452 then
	sram_write <= x"03DC0024";
end if;
if first_state_sram_input_id = 10453 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10454 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10455 then
	sram_write <= x"8200078C";
end if;
if first_state_sram_input_id = 10456 then
	sram_write <= x"07DC0024";
end if;
if first_state_sram_input_id = 10457 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 10458 then
	sram_write <= x"C05C000C";
end if;
if first_state_sram_input_id = 10459 then
	sram_write <= x"C07C0008";
end if;
if first_state_sram_input_id = 10460 then
	sram_write <= x"C09C0010";
end if;
if first_state_sram_input_id = 10461 then
	sram_write <= x"C0BC0004";
end if;
if first_state_sram_input_id = 10462 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10463 then
	sram_write <= x"03DC0024";
end if;
if first_state_sram_input_id = 10464 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10465 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10466 then
	sram_write <= x"82009C7C";
end if;
if first_state_sram_input_id = 10467 then
	sram_write <= x"07DC0024";
end if;
if first_state_sram_input_id = 10468 then
	sram_write <= x"C03C000C";
end if;
if first_state_sram_input_id = 10469 then
	sram_write <= x"02420001";
end if;
if first_state_sram_input_id = 10470 then
	sram_write <= x"C03C0000";
end if;
if first_state_sram_input_id = 10471 then
	sram_write <= x"02220002";
end if;
if first_state_sram_input_id = 10472 then
	sram_write <= x"02600005";
end if;
if first_state_sram_input_id = 10473 then
	sram_write <= x"8626A3B0";
end if;
if first_state_sram_input_id = 10474 then
	sram_write <= x"06620005";
end if;
if first_state_sram_input_id = 10475 then
	sram_write <= x"8200A3B4";
end if;
if first_state_sram_input_id = 10476 then
	sram_write <= x"00620000";
end if;
if first_state_sram_input_id = 10477 then
	sram_write <= x"C03C0014";
end if;
if first_state_sram_input_id = 10478 then
	sram_write <= x"C0820004";
end if;
if first_state_sram_input_id = 10479 then
	sram_write <= x"8648A3C4";
end if;
if first_state_sram_input_id = 10480 then
	sram_write <= x"8200A478";
end if;
if first_state_sram_input_id = 10481 then
	sram_write <= x"C0220004";
end if;
if first_state_sram_input_id = 10482 then
	sram_write <= x"06220001";
end if;
if first_state_sram_input_id = 10483 then
	sram_write <= x"C47C001C";
end if;
if first_state_sram_input_id = 10484 then
	sram_write <= x"C45C0020";
end if;
if first_state_sram_input_id = 10485 then
	sram_write <= x"8642A3DC";
end if;
if first_state_sram_input_id = 10486 then
	sram_write <= x"8200A404";
end if;
if first_state_sram_input_id = 10487 then
	sram_write <= x"02240001";
end if;
if first_state_sram_input_id = 10488 then
	sram_write <= x"C09C0008";
end if;
if first_state_sram_input_id = 10489 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10490 then
	sram_write <= x"00420000";
end if;
if first_state_sram_input_id = 10491 then
	sram_write <= x"00280000";
end if;
if first_state_sram_input_id = 10492 then
	sram_write <= x"03DC002C";
end if;
if first_state_sram_input_id = 10493 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10494 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10495 then
	sram_write <= x"82009C08";
end if;
if first_state_sram_input_id = 10496 then
	sram_write <= x"07DC002C";
end if;
if first_state_sram_input_id = 10497 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 10498 then
	sram_write <= x"C05C0020";
end if;
if first_state_sram_input_id = 10499 then
	sram_write <= x"C07C0010";
end if;
if first_state_sram_input_id = 10500 then
	sram_write <= x"C09C0004";
end if;
if first_state_sram_input_id = 10501 then
	sram_write <= x"C0BC0008";
end if;
if first_state_sram_input_id = 10502 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10503 then
	sram_write <= x"03DC002C";
end if;
if first_state_sram_input_id = 10504 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10505 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10506 then
	sram_write <= x"82009C7C";
end if;
if first_state_sram_input_id = 10507 then
	sram_write <= x"07DC002C";
end if;
if first_state_sram_input_id = 10508 then
	sram_write <= x"C03C0020";
end if;
if first_state_sram_input_id = 10509 then
	sram_write <= x"02220001";
end if;
if first_state_sram_input_id = 10510 then
	sram_write <= x"C05C001C";
end if;
if first_state_sram_input_id = 10511 then
	sram_write <= x"02440002";
end if;
if first_state_sram_input_id = 10512 then
	sram_write <= x"02600005";
end if;
if first_state_sram_input_id = 10513 then
	sram_write <= x"8646A450";
end if;
if first_state_sram_input_id = 10514 then
	sram_write <= x"06A40005";
end if;
if first_state_sram_input_id = 10515 then
	sram_write <= x"8200A454";
end if;
if first_state_sram_input_id = 10516 then
	sram_write <= x"00A40000";
end if;
if first_state_sram_input_id = 10517 then
	sram_write <= x"C05C0004";
end if;
if first_state_sram_input_id = 10518 then
	sram_write <= x"C07C0008";
end if;
if first_state_sram_input_id = 10519 then
	sram_write <= x"C09C0010";
end if;
if first_state_sram_input_id = 10520 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10521 then
	sram_write <= x"03DC002C";
end if;
if first_state_sram_input_id = 10522 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10523 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10524 then
	sram_write <= x"8200A164";
end if;
if first_state_sram_input_id = 10525 then
	sram_write <= x"07DC002C";
end if;
if first_state_sram_input_id = 10526 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 10527 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 10528 then
	sram_write <= x"40200000";
end if;
if first_state_sram_input_id = 10529 then
	sram_write <= x"CC3C0000";
end if;
if first_state_sram_input_id = 10530 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10531 then
	sram_write <= x"03DC0010";
end if;
if first_state_sram_input_id = 10532 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10533 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10534 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 10535 then
	sram_write <= x"07DC0010";
end if;
if first_state_sram_input_id = 10536 then
	sram_write <= x"02400003";
end if;
if first_state_sram_input_id = 10537 then
	sram_write <= x"C83C0000";
end if;
if first_state_sram_input_id = 10538 then
	sram_write <= x"C43C0008";
end if;
if first_state_sram_input_id = 10539 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10540 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 10541 then
	sram_write <= x"03DC0014";
end if;
if first_state_sram_input_id = 10542 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10543 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10544 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 10545 then
	sram_write <= x"07DC0014";
end if;
if first_state_sram_input_id = 10546 then
	sram_write <= x"00420000";
end if;
if first_state_sram_input_id = 10547 then
	sram_write <= x"02200005";
end if;
if first_state_sram_input_id = 10548 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10549 then
	sram_write <= x"03DC0014";
end if;
if first_state_sram_input_id = 10550 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10551 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10552 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 10553 then
	sram_write <= x"07DC0014";
end if;
if first_state_sram_input_id = 10554 then
	sram_write <= x"02400003";
end if;
if first_state_sram_input_id = 10555 then
	sram_write <= x"C83C0000";
end if;
if first_state_sram_input_id = 10556 then
	sram_write <= x"C43C000C";
end if;
if first_state_sram_input_id = 10557 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10558 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 10559 then
	sram_write <= x"03DC0018";
end if;
if first_state_sram_input_id = 10560 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10561 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10562 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 10563 then
	sram_write <= x"07DC0018";
end if;
if first_state_sram_input_id = 10564 then
	sram_write <= x"C05C000C";
end if;
if first_state_sram_input_id = 10565 then
	sram_write <= x"C4240004";
end if;
if first_state_sram_input_id = 10566 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 10567 then
	sram_write <= x"C83C0000";
end if;
if first_state_sram_input_id = 10568 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10569 then
	sram_write <= x"03DC0018";
end if;
if first_state_sram_input_id = 10570 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10571 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10572 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 10573 then
	sram_write <= x"07DC0018";
end if;
if first_state_sram_input_id = 10574 then
	sram_write <= x"C05C000C";
end if;
if first_state_sram_input_id = 10575 then
	sram_write <= x"C4240008";
end if;
if first_state_sram_input_id = 10576 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 10577 then
	sram_write <= x"C83C0000";
end if;
if first_state_sram_input_id = 10578 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10579 then
	sram_write <= x"03DC0018";
end if;
if first_state_sram_input_id = 10580 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10581 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10582 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 10583 then
	sram_write <= x"07DC0018";
end if;
if first_state_sram_input_id = 10584 then
	sram_write <= x"C05C000C";
end if;
if first_state_sram_input_id = 10585 then
	sram_write <= x"C424000C";
end if;
if first_state_sram_input_id = 10586 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 10587 then
	sram_write <= x"C83C0000";
end if;
if first_state_sram_input_id = 10588 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10589 then
	sram_write <= x"03DC0018";
end if;
if first_state_sram_input_id = 10590 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10591 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10592 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 10593 then
	sram_write <= x"07DC0018";
end if;
if first_state_sram_input_id = 10594 then
	sram_write <= x"C05C000C";
end if;
if first_state_sram_input_id = 10595 then
	sram_write <= x"C4240010";
end if;
if first_state_sram_input_id = 10596 then
	sram_write <= x"02200005";
end if;
if first_state_sram_input_id = 10597 then
	sram_write <= x"02600000";
end if;
if first_state_sram_input_id = 10598 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10599 then
	sram_write <= x"00460000";
end if;
if first_state_sram_input_id = 10600 then
	sram_write <= x"03DC0018";
end if;
if first_state_sram_input_id = 10601 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10602 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10603 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 10604 then
	sram_write <= x"07DC0018";
end if;
if first_state_sram_input_id = 10605 then
	sram_write <= x"02400005";
end if;
if first_state_sram_input_id = 10606 then
	sram_write <= x"02600000";
end if;
if first_state_sram_input_id = 10607 then
	sram_write <= x"C43C0010";
end if;
if first_state_sram_input_id = 10608 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10609 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 10610 then
	sram_write <= x"00460000";
end if;
if first_state_sram_input_id = 10611 then
	sram_write <= x"03DC001C";
end if;
if first_state_sram_input_id = 10612 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10613 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10614 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 10615 then
	sram_write <= x"07DC001C";
end if;
if first_state_sram_input_id = 10616 then
	sram_write <= x"02400003";
end if;
if first_state_sram_input_id = 10617 then
	sram_write <= x"C83C0000";
end if;
if first_state_sram_input_id = 10618 then
	sram_write <= x"C43C0014";
end if;
if first_state_sram_input_id = 10619 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10620 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 10621 then
	sram_write <= x"03DC0020";
end if;
if first_state_sram_input_id = 10622 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10623 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10624 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 10625 then
	sram_write <= x"07DC0020";
end if;
if first_state_sram_input_id = 10626 then
	sram_write <= x"00420000";
end if;
if first_state_sram_input_id = 10627 then
	sram_write <= x"02200005";
end if;
if first_state_sram_input_id = 10628 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10629 then
	sram_write <= x"03DC0020";
end if;
if first_state_sram_input_id = 10630 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10631 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10632 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 10633 then
	sram_write <= x"07DC0020";
end if;
if first_state_sram_input_id = 10634 then
	sram_write <= x"02400003";
end if;
if first_state_sram_input_id = 10635 then
	sram_write <= x"C83C0000";
end if;
if first_state_sram_input_id = 10636 then
	sram_write <= x"C43C0018";
end if;
if first_state_sram_input_id = 10637 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10638 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 10639 then
	sram_write <= x"03DC0024";
end if;
if first_state_sram_input_id = 10640 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10641 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10642 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 10643 then
	sram_write <= x"07DC0024";
end if;
if first_state_sram_input_id = 10644 then
	sram_write <= x"C05C0018";
end if;
if first_state_sram_input_id = 10645 then
	sram_write <= x"C4240004";
end if;
if first_state_sram_input_id = 10646 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 10647 then
	sram_write <= x"C83C0000";
end if;
if first_state_sram_input_id = 10648 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10649 then
	sram_write <= x"03DC0024";
end if;
if first_state_sram_input_id = 10650 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10651 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10652 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 10653 then
	sram_write <= x"07DC0024";
end if;
if first_state_sram_input_id = 10654 then
	sram_write <= x"C05C0018";
end if;
if first_state_sram_input_id = 10655 then
	sram_write <= x"C4240008";
end if;
if first_state_sram_input_id = 10656 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 10657 then
	sram_write <= x"C83C0000";
end if;
if first_state_sram_input_id = 10658 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10659 then
	sram_write <= x"03DC0024";
end if;
if first_state_sram_input_id = 10660 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10661 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10662 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 10663 then
	sram_write <= x"07DC0024";
end if;
if first_state_sram_input_id = 10664 then
	sram_write <= x"C05C0018";
end if;
if first_state_sram_input_id = 10665 then
	sram_write <= x"C424000C";
end if;
if first_state_sram_input_id = 10666 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 10667 then
	sram_write <= x"C83C0000";
end if;
if first_state_sram_input_id = 10668 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10669 then
	sram_write <= x"03DC0024";
end if;
if first_state_sram_input_id = 10670 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10671 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10672 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 10673 then
	sram_write <= x"07DC0024";
end if;
if first_state_sram_input_id = 10674 then
	sram_write <= x"C05C0018";
end if;
if first_state_sram_input_id = 10675 then
	sram_write <= x"C4240010";
end if;
if first_state_sram_input_id = 10676 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 10677 then
	sram_write <= x"C83C0000";
end if;
if first_state_sram_input_id = 10678 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10679 then
	sram_write <= x"03DC0024";
end if;
if first_state_sram_input_id = 10680 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10681 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10682 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 10683 then
	sram_write <= x"07DC0024";
end if;
if first_state_sram_input_id = 10684 then
	sram_write <= x"00420000";
end if;
if first_state_sram_input_id = 10685 then
	sram_write <= x"02200005";
end if;
if first_state_sram_input_id = 10686 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10687 then
	sram_write <= x"03DC0024";
end if;
if first_state_sram_input_id = 10688 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10689 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10690 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 10691 then
	sram_write <= x"07DC0024";
end if;
if first_state_sram_input_id = 10692 then
	sram_write <= x"02400003";
end if;
if first_state_sram_input_id = 10693 then
	sram_write <= x"C83C0000";
end if;
if first_state_sram_input_id = 10694 then
	sram_write <= x"C43C001C";
end if;
if first_state_sram_input_id = 10695 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10696 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 10697 then
	sram_write <= x"03DC0028";
end if;
if first_state_sram_input_id = 10698 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10699 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10700 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 10701 then
	sram_write <= x"07DC0028";
end if;
if first_state_sram_input_id = 10702 then
	sram_write <= x"C05C001C";
end if;
if first_state_sram_input_id = 10703 then
	sram_write <= x"C4240004";
end if;
if first_state_sram_input_id = 10704 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 10705 then
	sram_write <= x"C83C0000";
end if;
if first_state_sram_input_id = 10706 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10707 then
	sram_write <= x"03DC0028";
end if;
if first_state_sram_input_id = 10708 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10709 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10710 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 10711 then
	sram_write <= x"07DC0028";
end if;
if first_state_sram_input_id = 10712 then
	sram_write <= x"C05C001C";
end if;
if first_state_sram_input_id = 10713 then
	sram_write <= x"C4240008";
end if;
if first_state_sram_input_id = 10714 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 10715 then
	sram_write <= x"C83C0000";
end if;
if first_state_sram_input_id = 10716 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10717 then
	sram_write <= x"03DC0028";
end if;
if first_state_sram_input_id = 10718 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10719 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10720 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 10721 then
	sram_write <= x"07DC0028";
end if;
if first_state_sram_input_id = 10722 then
	sram_write <= x"C05C001C";
end if;
if first_state_sram_input_id = 10723 then
	sram_write <= x"C424000C";
end if;
if first_state_sram_input_id = 10724 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 10725 then
	sram_write <= x"C83C0000";
end if;
if first_state_sram_input_id = 10726 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10727 then
	sram_write <= x"03DC0028";
end if;
if first_state_sram_input_id = 10728 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10729 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10730 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 10731 then
	sram_write <= x"07DC0028";
end if;
if first_state_sram_input_id = 10732 then
	sram_write <= x"C05C001C";
end if;
if first_state_sram_input_id = 10733 then
	sram_write <= x"C4240010";
end if;
if first_state_sram_input_id = 10734 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 10735 then
	sram_write <= x"02600000";
end if;
if first_state_sram_input_id = 10736 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10737 then
	sram_write <= x"00460000";
end if;
if first_state_sram_input_id = 10738 then
	sram_write <= x"03DC0028";
end if;
if first_state_sram_input_id = 10739 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10740 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10741 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 10742 then
	sram_write <= x"07DC0028";
end if;
if first_state_sram_input_id = 10743 then
	sram_write <= x"02400003";
end if;
if first_state_sram_input_id = 10744 then
	sram_write <= x"C83C0000";
end if;
if first_state_sram_input_id = 10745 then
	sram_write <= x"C43C0020";
end if;
if first_state_sram_input_id = 10746 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10747 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 10748 then
	sram_write <= x"03DC002C";
end if;
if first_state_sram_input_id = 10749 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10750 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10751 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 10752 then
	sram_write <= x"07DC002C";
end if;
if first_state_sram_input_id = 10753 then
	sram_write <= x"00420000";
end if;
if first_state_sram_input_id = 10754 then
	sram_write <= x"02200005";
end if;
if first_state_sram_input_id = 10755 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10756 then
	sram_write <= x"03DC002C";
end if;
if first_state_sram_input_id = 10757 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10758 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10759 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 10760 then
	sram_write <= x"07DC002C";
end if;
if first_state_sram_input_id = 10761 then
	sram_write <= x"02400003";
end if;
if first_state_sram_input_id = 10762 then
	sram_write <= x"C83C0000";
end if;
if first_state_sram_input_id = 10763 then
	sram_write <= x"C43C0024";
end if;
if first_state_sram_input_id = 10764 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10765 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 10766 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 10767 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10768 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10769 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 10770 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 10771 then
	sram_write <= x"C05C0024";
end if;
if first_state_sram_input_id = 10772 then
	sram_write <= x"C4240004";
end if;
if first_state_sram_input_id = 10773 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 10774 then
	sram_write <= x"C83C0000";
end if;
if first_state_sram_input_id = 10775 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10776 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 10777 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10778 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10779 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 10780 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 10781 then
	sram_write <= x"C05C0024";
end if;
if first_state_sram_input_id = 10782 then
	sram_write <= x"C4240008";
end if;
if first_state_sram_input_id = 10783 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 10784 then
	sram_write <= x"C83C0000";
end if;
if first_state_sram_input_id = 10785 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10786 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 10787 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10788 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10789 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 10790 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 10791 then
	sram_write <= x"C05C0024";
end if;
if first_state_sram_input_id = 10792 then
	sram_write <= x"C424000C";
end if;
if first_state_sram_input_id = 10793 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 10794 then
	sram_write <= x"C83C0000";
end if;
if first_state_sram_input_id = 10795 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10796 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 10797 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10798 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10799 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 10800 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 10801 then
	sram_write <= x"C05C0024";
end if;
if first_state_sram_input_id = 10802 then
	sram_write <= x"C4240010";
end if;
if first_state_sram_input_id = 10803 then
	sram_write <= x"003A0000";
end if;
if first_state_sram_input_id = 10804 then
	sram_write <= x"03BA0020";
end if;
if first_state_sram_input_id = 10805 then
	sram_write <= x"C442001C";
end if;
if first_state_sram_input_id = 10806 then
	sram_write <= x"C05C0020";
end if;
if first_state_sram_input_id = 10807 then
	sram_write <= x"C4420018";
end if;
if first_state_sram_input_id = 10808 then
	sram_write <= x"C05C001C";
end if;
if first_state_sram_input_id = 10809 then
	sram_write <= x"C4420014";
end if;
if first_state_sram_input_id = 10810 then
	sram_write <= x"C05C0018";
end if;
if first_state_sram_input_id = 10811 then
	sram_write <= x"C4420010";
end if;
if first_state_sram_input_id = 10812 then
	sram_write <= x"C05C0014";
end if;
if first_state_sram_input_id = 10813 then
	sram_write <= x"C442000C";
end if;
if first_state_sram_input_id = 10814 then
	sram_write <= x"C05C0010";
end if;
if first_state_sram_input_id = 10815 then
	sram_write <= x"C4420008";
end if;
if first_state_sram_input_id = 10816 then
	sram_write <= x"C05C000C";
end if;
if first_state_sram_input_id = 10817 then
	sram_write <= x"C4420004";
end if;
if first_state_sram_input_id = 10818 then
	sram_write <= x"C05C0008";
end if;
if first_state_sram_input_id = 10819 then
	sram_write <= x"C4420000";
end if;
if first_state_sram_input_id = 10820 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 10821 then
	sram_write <= x"8640AE10";
end if;
if first_state_sram_input_id = 10822 then
	sram_write <= x"02600003";
end if;
if first_state_sram_input_id = 10823 then
	sram_write <= x"40200000";
end if;
if first_state_sram_input_id = 10824 then
	sram_write <= x"C43C0000";
end if;
if first_state_sram_input_id = 10825 then
	sram_write <= x"C45C0004";
end if;
if first_state_sram_input_id = 10826 then
	sram_write <= x"CC3C0008";
end if;
if first_state_sram_input_id = 10827 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10828 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 10829 then
	sram_write <= x"03DC0018";
end if;
if first_state_sram_input_id = 10830 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10831 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10832 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 10833 then
	sram_write <= x"07DC0018";
end if;
if first_state_sram_input_id = 10834 then
	sram_write <= x"02400003";
end if;
if first_state_sram_input_id = 10835 then
	sram_write <= x"C83C0008";
end if;
if first_state_sram_input_id = 10836 then
	sram_write <= x"C43C0010";
end if;
if first_state_sram_input_id = 10837 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10838 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 10839 then
	sram_write <= x"03DC001C";
end if;
if first_state_sram_input_id = 10840 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10841 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10842 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 10843 then
	sram_write <= x"07DC001C";
end if;
if first_state_sram_input_id = 10844 then
	sram_write <= x"00420000";
end if;
if first_state_sram_input_id = 10845 then
	sram_write <= x"02200005";
end if;
if first_state_sram_input_id = 10846 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10847 then
	sram_write <= x"03DC001C";
end if;
if first_state_sram_input_id = 10848 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10849 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10850 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 10851 then
	sram_write <= x"07DC001C";
end if;
if first_state_sram_input_id = 10852 then
	sram_write <= x"02400003";
end if;
if first_state_sram_input_id = 10853 then
	sram_write <= x"C83C0008";
end if;
if first_state_sram_input_id = 10854 then
	sram_write <= x"C43C0014";
end if;
if first_state_sram_input_id = 10855 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10856 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 10857 then
	sram_write <= x"03DC0020";
end if;
if first_state_sram_input_id = 10858 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10859 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10860 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 10861 then
	sram_write <= x"07DC0020";
end if;
if first_state_sram_input_id = 10862 then
	sram_write <= x"C05C0014";
end if;
if first_state_sram_input_id = 10863 then
	sram_write <= x"C4240004";
end if;
if first_state_sram_input_id = 10864 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 10865 then
	sram_write <= x"C83C0008";
end if;
if first_state_sram_input_id = 10866 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10867 then
	sram_write <= x"03DC0020";
end if;
if first_state_sram_input_id = 10868 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10869 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10870 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 10871 then
	sram_write <= x"07DC0020";
end if;
if first_state_sram_input_id = 10872 then
	sram_write <= x"C05C0014";
end if;
if first_state_sram_input_id = 10873 then
	sram_write <= x"C4240008";
end if;
if first_state_sram_input_id = 10874 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 10875 then
	sram_write <= x"C83C0008";
end if;
if first_state_sram_input_id = 10876 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10877 then
	sram_write <= x"03DC0020";
end if;
if first_state_sram_input_id = 10878 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10879 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10880 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 10881 then
	sram_write <= x"07DC0020";
end if;
if first_state_sram_input_id = 10882 then
	sram_write <= x"C05C0014";
end if;
if first_state_sram_input_id = 10883 then
	sram_write <= x"C424000C";
end if;
if first_state_sram_input_id = 10884 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 10885 then
	sram_write <= x"C83C0008";
end if;
if first_state_sram_input_id = 10886 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10887 then
	sram_write <= x"03DC0020";
end if;
if first_state_sram_input_id = 10888 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10889 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10890 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 10891 then
	sram_write <= x"07DC0020";
end if;
if first_state_sram_input_id = 10892 then
	sram_write <= x"C05C0014";
end if;
if first_state_sram_input_id = 10893 then
	sram_write <= x"C4240010";
end if;
if first_state_sram_input_id = 10894 then
	sram_write <= x"02200005";
end if;
if first_state_sram_input_id = 10895 then
	sram_write <= x"02600000";
end if;
if first_state_sram_input_id = 10896 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10897 then
	sram_write <= x"00460000";
end if;
if first_state_sram_input_id = 10898 then
	sram_write <= x"03DC0020";
end if;
if first_state_sram_input_id = 10899 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10900 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10901 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 10902 then
	sram_write <= x"07DC0020";
end if;
if first_state_sram_input_id = 10903 then
	sram_write <= x"02400005";
end if;
if first_state_sram_input_id = 10904 then
	sram_write <= x"02600000";
end if;
if first_state_sram_input_id = 10905 then
	sram_write <= x"C43C0018";
end if;
if first_state_sram_input_id = 10906 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10907 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 10908 then
	sram_write <= x"00460000";
end if;
if first_state_sram_input_id = 10909 then
	sram_write <= x"03DC0024";
end if;
if first_state_sram_input_id = 10910 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10911 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10912 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 10913 then
	sram_write <= x"07DC0024";
end if;
if first_state_sram_input_id = 10914 then
	sram_write <= x"02400003";
end if;
if first_state_sram_input_id = 10915 then
	sram_write <= x"C83C0008";
end if;
if first_state_sram_input_id = 10916 then
	sram_write <= x"C43C001C";
end if;
if first_state_sram_input_id = 10917 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10918 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 10919 then
	sram_write <= x"03DC0028";
end if;
if first_state_sram_input_id = 10920 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10921 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10922 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 10923 then
	sram_write <= x"07DC0028";
end if;
if first_state_sram_input_id = 10924 then
	sram_write <= x"00420000";
end if;
if first_state_sram_input_id = 10925 then
	sram_write <= x"02200005";
end if;
if first_state_sram_input_id = 10926 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10927 then
	sram_write <= x"03DC0028";
end if;
if first_state_sram_input_id = 10928 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10929 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10930 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 10931 then
	sram_write <= x"07DC0028";
end if;
if first_state_sram_input_id = 10932 then
	sram_write <= x"02400003";
end if;
if first_state_sram_input_id = 10933 then
	sram_write <= x"C83C0008";
end if;
if first_state_sram_input_id = 10934 then
	sram_write <= x"C43C0020";
end if;
if first_state_sram_input_id = 10935 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10936 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 10937 then
	sram_write <= x"03DC002C";
end if;
if first_state_sram_input_id = 10938 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10939 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10940 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 10941 then
	sram_write <= x"07DC002C";
end if;
if first_state_sram_input_id = 10942 then
	sram_write <= x"C05C0020";
end if;
if first_state_sram_input_id = 10943 then
	sram_write <= x"C4240004";
end if;
if first_state_sram_input_id = 10944 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 10945 then
	sram_write <= x"C83C0008";
end if;
if first_state_sram_input_id = 10946 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10947 then
	sram_write <= x"03DC002C";
end if;
if first_state_sram_input_id = 10948 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10949 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10950 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 10951 then
	sram_write <= x"07DC002C";
end if;
if first_state_sram_input_id = 10952 then
	sram_write <= x"C05C0020";
end if;
if first_state_sram_input_id = 10953 then
	sram_write <= x"C4240008";
end if;
if first_state_sram_input_id = 10954 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 10955 then
	sram_write <= x"C83C0008";
end if;
if first_state_sram_input_id = 10956 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10957 then
	sram_write <= x"03DC002C";
end if;
if first_state_sram_input_id = 10958 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10959 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10960 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 10961 then
	sram_write <= x"07DC002C";
end if;
if first_state_sram_input_id = 10962 then
	sram_write <= x"C05C0020";
end if;
if first_state_sram_input_id = 10963 then
	sram_write <= x"C424000C";
end if;
if first_state_sram_input_id = 10964 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 10965 then
	sram_write <= x"C83C0008";
end if;
if first_state_sram_input_id = 10966 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10967 then
	sram_write <= x"03DC002C";
end if;
if first_state_sram_input_id = 10968 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10969 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10970 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 10971 then
	sram_write <= x"07DC002C";
end if;
if first_state_sram_input_id = 10972 then
	sram_write <= x"C05C0020";
end if;
if first_state_sram_input_id = 10973 then
	sram_write <= x"C4240010";
end if;
if first_state_sram_input_id = 10974 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 10975 then
	sram_write <= x"C83C0008";
end if;
if first_state_sram_input_id = 10976 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10977 then
	sram_write <= x"03DC002C";
end if;
if first_state_sram_input_id = 10978 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10979 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10980 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 10981 then
	sram_write <= x"07DC002C";
end if;
if first_state_sram_input_id = 10982 then
	sram_write <= x"00420000";
end if;
if first_state_sram_input_id = 10983 then
	sram_write <= x"02200005";
end if;
if first_state_sram_input_id = 10984 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10985 then
	sram_write <= x"03DC002C";
end if;
if first_state_sram_input_id = 10986 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10987 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10988 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 10989 then
	sram_write <= x"07DC002C";
end if;
if first_state_sram_input_id = 10990 then
	sram_write <= x"02400003";
end if;
if first_state_sram_input_id = 10991 then
	sram_write <= x"C83C0008";
end if;
if first_state_sram_input_id = 10992 then
	sram_write <= x"C43C0024";
end if;
if first_state_sram_input_id = 10993 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 10994 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 10995 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 10996 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 10997 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 10998 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 10999 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 11000 then
	sram_write <= x"C05C0024";
end if;
if first_state_sram_input_id = 11001 then
	sram_write <= x"C4240004";
end if;
if first_state_sram_input_id = 11002 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 11003 then
	sram_write <= x"C83C0008";
end if;
if first_state_sram_input_id = 11004 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11005 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 11006 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11007 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11008 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 11009 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 11010 then
	sram_write <= x"C05C0024";
end if;
if first_state_sram_input_id = 11011 then
	sram_write <= x"C4240008";
end if;
if first_state_sram_input_id = 11012 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 11013 then
	sram_write <= x"C83C0008";
end if;
if first_state_sram_input_id = 11014 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11015 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 11016 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11017 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11018 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 11019 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 11020 then
	sram_write <= x"C05C0024";
end if;
if first_state_sram_input_id = 11021 then
	sram_write <= x"C424000C";
end if;
if first_state_sram_input_id = 11022 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 11023 then
	sram_write <= x"C83C0008";
end if;
if first_state_sram_input_id = 11024 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11025 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 11026 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11027 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11028 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 11029 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 11030 then
	sram_write <= x"C05C0024";
end if;
if first_state_sram_input_id = 11031 then
	sram_write <= x"C4240010";
end if;
if first_state_sram_input_id = 11032 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 11033 then
	sram_write <= x"02600000";
end if;
if first_state_sram_input_id = 11034 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11035 then
	sram_write <= x"00460000";
end if;
if first_state_sram_input_id = 11036 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 11037 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11038 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11039 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 11040 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 11041 then
	sram_write <= x"02400003";
end if;
if first_state_sram_input_id = 11042 then
	sram_write <= x"C83C0008";
end if;
if first_state_sram_input_id = 11043 then
	sram_write <= x"C43C0028";
end if;
if first_state_sram_input_id = 11044 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11045 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 11046 then
	sram_write <= x"03DC0034";
end if;
if first_state_sram_input_id = 11047 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11048 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11049 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 11050 then
	sram_write <= x"07DC0034";
end if;
if first_state_sram_input_id = 11051 then
	sram_write <= x"00420000";
end if;
if first_state_sram_input_id = 11052 then
	sram_write <= x"02200005";
end if;
if first_state_sram_input_id = 11053 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11054 then
	sram_write <= x"03DC0034";
end if;
if first_state_sram_input_id = 11055 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11056 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11057 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 11058 then
	sram_write <= x"07DC0034";
end if;
if first_state_sram_input_id = 11059 then
	sram_write <= x"02400003";
end if;
if first_state_sram_input_id = 11060 then
	sram_write <= x"C83C0008";
end if;
if first_state_sram_input_id = 11061 then
	sram_write <= x"C43C002C";
end if;
if first_state_sram_input_id = 11062 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11063 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 11064 then
	sram_write <= x"03DC0038";
end if;
if first_state_sram_input_id = 11065 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11066 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11067 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 11068 then
	sram_write <= x"07DC0038";
end if;
if first_state_sram_input_id = 11069 then
	sram_write <= x"C05C002C";
end if;
if first_state_sram_input_id = 11070 then
	sram_write <= x"C4240004";
end if;
if first_state_sram_input_id = 11071 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 11072 then
	sram_write <= x"C83C0008";
end if;
if first_state_sram_input_id = 11073 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11074 then
	sram_write <= x"03DC0038";
end if;
if first_state_sram_input_id = 11075 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11076 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11077 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 11078 then
	sram_write <= x"07DC0038";
end if;
if first_state_sram_input_id = 11079 then
	sram_write <= x"C05C002C";
end if;
if first_state_sram_input_id = 11080 then
	sram_write <= x"C4240008";
end if;
if first_state_sram_input_id = 11081 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 11082 then
	sram_write <= x"C83C0008";
end if;
if first_state_sram_input_id = 11083 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11084 then
	sram_write <= x"03DC0038";
end if;
if first_state_sram_input_id = 11085 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11086 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11087 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 11088 then
	sram_write <= x"07DC0038";
end if;
if first_state_sram_input_id = 11089 then
	sram_write <= x"C05C002C";
end if;
if first_state_sram_input_id = 11090 then
	sram_write <= x"C424000C";
end if;
if first_state_sram_input_id = 11091 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 11092 then
	sram_write <= x"C83C0008";
end if;
if first_state_sram_input_id = 11093 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11094 then
	sram_write <= x"03DC0038";
end if;
if first_state_sram_input_id = 11095 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11096 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11097 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 11098 then
	sram_write <= x"07DC0038";
end if;
if first_state_sram_input_id = 11099 then
	sram_write <= x"C05C002C";
end if;
if first_state_sram_input_id = 11100 then
	sram_write <= x"C4240010";
end if;
if first_state_sram_input_id = 11101 then
	sram_write <= x"003A0000";
end if;
if first_state_sram_input_id = 11102 then
	sram_write <= x"03BA0020";
end if;
if first_state_sram_input_id = 11103 then
	sram_write <= x"C442001C";
end if;
if first_state_sram_input_id = 11104 then
	sram_write <= x"C05C0028";
end if;
if first_state_sram_input_id = 11105 then
	sram_write <= x"C4420018";
end if;
if first_state_sram_input_id = 11106 then
	sram_write <= x"C05C0024";
end if;
if first_state_sram_input_id = 11107 then
	sram_write <= x"C4420014";
end if;
if first_state_sram_input_id = 11108 then
	sram_write <= x"C05C0020";
end if;
if first_state_sram_input_id = 11109 then
	sram_write <= x"C4420010";
end if;
if first_state_sram_input_id = 11110 then
	sram_write <= x"C05C001C";
end if;
if first_state_sram_input_id = 11111 then
	sram_write <= x"C442000C";
end if;
if first_state_sram_input_id = 11112 then
	sram_write <= x"C05C0018";
end if;
if first_state_sram_input_id = 11113 then
	sram_write <= x"C4420008";
end if;
if first_state_sram_input_id = 11114 then
	sram_write <= x"C05C0014";
end if;
if first_state_sram_input_id = 11115 then
	sram_write <= x"C4420004";
end if;
if first_state_sram_input_id = 11116 then
	sram_write <= x"C05C0010";
end if;
if first_state_sram_input_id = 11117 then
	sram_write <= x"C4420000";
end if;
if first_state_sram_input_id = 11118 then
	sram_write <= x"C05C0004";
end if;
if first_state_sram_input_id = 11119 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 11120 then
	sram_write <= x"C09C0000";
end if;
if first_state_sram_input_id = 11121 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 11122 then
	sram_write <= x"06240001";
end if;
if first_state_sram_input_id = 11123 then
	sram_write <= x"8620AE08";
end if;
if first_state_sram_input_id = 11124 then
	sram_write <= x"C43C0030";
end if;
if first_state_sram_input_id = 11125 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11126 then
	sram_write <= x"03DC003C";
end if;
if first_state_sram_input_id = 11127 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11128 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11129 then
	sram_write <= x"8200A47C";
end if;
if first_state_sram_input_id = 11130 then
	sram_write <= x"07DC003C";
end if;
if first_state_sram_input_id = 11131 then
	sram_write <= x"C05C0030";
end if;
if first_state_sram_input_id = 11132 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 11133 then
	sram_write <= x"C09C0000";
end if;
if first_state_sram_input_id = 11134 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 11135 then
	sram_write <= x"06440001";
end if;
if first_state_sram_input_id = 11136 then
	sram_write <= x"00280000";
end if;
if first_state_sram_input_id = 11137 then
	sram_write <= x"8200A914";
end if;
if first_state_sram_input_id = 11138 then
	sram_write <= x"00280000";
end if;
if first_state_sram_input_id = 11139 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 11140 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 11141 then
	sram_write <= x"02800005";
end if;
if first_state_sram_input_id = 11142 then
	sram_write <= x"8628AFA0";
end if;
if first_state_sram_input_id = 11143 then
	sram_write <= x"48622000";
end if;
if first_state_sram_input_id = 11144 then
	sram_write <= x"48844000";
end if;
if first_state_sram_input_id = 11145 then
	sram_write <= x"40668000";
end if;
if first_state_sram_input_id = 11146 then
	sram_write <= x"C88000A8";
end if;
if first_state_sram_input_id = 11147 then
	sram_write <= x"40668000";
end if;
if first_state_sram_input_id = 11148 then
	sram_write <= x"C47C0000";
end if;
if first_state_sram_input_id = 11149 then
	sram_write <= x"C45C0004";
end if;
if first_state_sram_input_id = 11150 then
	sram_write <= x"CC5C0008";
end if;
if first_state_sram_input_id = 11151 then
	sram_write <= x"CC3C0010";
end if;
if first_state_sram_input_id = 11152 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11153 then
	sram_write <= x"40206000";
end if;
if first_state_sram_input_id = 11154 then
	sram_write <= x"03DC0020";
end if;
if first_state_sram_input_id = 11155 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11156 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11157 then
	sram_write <= x"8200083C";
end if;
if first_state_sram_input_id = 11158 then
	sram_write <= x"07DC0020";
end if;
if first_state_sram_input_id = 11159 then
	sram_write <= x"CC3C0018";
end if;
if first_state_sram_input_id = 11160 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11161 then
	sram_write <= x"03DC0028";
end if;
if first_state_sram_input_id = 11162 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11163 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11164 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 11165 then
	sram_write <= x"07DC0028";
end if;
if first_state_sram_input_id = 11166 then
	sram_write <= x"C85C0010";
end if;
if first_state_sram_input_id = 11167 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 11168 then
	sram_write <= x"C85C0018";
end if;
if first_state_sram_input_id = 11169 then
	sram_write <= x"CC3C0020";
end if;
if first_state_sram_input_id = 11170 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11171 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 11172 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 11173 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11174 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11175 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 11176 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 11177 then
	sram_write <= x"C85C0008";
end if;
if first_state_sram_input_id = 11178 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 11179 then
	sram_write <= x"C85C0018";
end if;
if first_state_sram_input_id = 11180 then
	sram_write <= x"CC3C0028";
end if;
if first_state_sram_input_id = 11181 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11182 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 11183 then
	sram_write <= x"03DC0038";
end if;
if first_state_sram_input_id = 11184 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11185 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11186 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 11187 then
	sram_write <= x"07DC0038";
end if;
if first_state_sram_input_id = 11188 then
	sram_write <= x"02200354";
end if;
if first_state_sram_input_id = 11189 then
	sram_write <= x"C05C0004";
end if;
if first_state_sram_input_id = 11190 then
	sram_write <= x"22440220";
end if;
if first_state_sram_input_id = 11191 then
	sram_write <= x"D0224000";
end if;
if first_state_sram_input_id = 11192 then
	sram_write <= x"C05C0000";
end if;
if first_state_sram_input_id = 11193 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 11194 then
	sram_write <= x"D0626000";
end if;
if first_state_sram_input_id = 11195 then
	sram_write <= x"C0660000";
end if;
if first_state_sram_input_id = 11196 then
	sram_write <= x"C85C0020";
end if;
if first_state_sram_input_id = 11197 then
	sram_write <= x"CC460000";
end if;
if first_state_sram_input_id = 11198 then
	sram_write <= x"C87C0028";
end if;
if first_state_sram_input_id = 11199 then
	sram_write <= x"CC660004";
end if;
if first_state_sram_input_id = 11200 then
	sram_write <= x"CC260008";
end if;
if first_state_sram_input_id = 11201 then
	sram_write <= x"02640028";
end if;
if first_state_sram_input_id = 11202 then
	sram_write <= x"22660220";
end if;
if first_state_sram_input_id = 11203 then
	sram_write <= x"D0626000";
end if;
if first_state_sram_input_id = 11204 then
	sram_write <= x"C0660000";
end if;
if first_state_sram_input_id = 11205 then
	sram_write <= x"44806000";
end if;
if first_state_sram_input_id = 11206 then
	sram_write <= x"CC460000";
end if;
if first_state_sram_input_id = 11207 then
	sram_write <= x"CC260004";
end if;
if first_state_sram_input_id = 11208 then
	sram_write <= x"CC860008";
end if;
if first_state_sram_input_id = 11209 then
	sram_write <= x"02640050";
end if;
if first_state_sram_input_id = 11210 then
	sram_write <= x"22660220";
end if;
if first_state_sram_input_id = 11211 then
	sram_write <= x"D0626000";
end if;
if first_state_sram_input_id = 11212 then
	sram_write <= x"C0660000";
end if;
if first_state_sram_input_id = 11213 then
	sram_write <= x"44A04000";
end if;
if first_state_sram_input_id = 11214 then
	sram_write <= x"CC260000";
end if;
if first_state_sram_input_id = 11215 then
	sram_write <= x"CCA60004";
end if;
if first_state_sram_input_id = 11216 then
	sram_write <= x"CC860008";
end if;
if first_state_sram_input_id = 11217 then
	sram_write <= x"02640001";
end if;
if first_state_sram_input_id = 11218 then
	sram_write <= x"22660220";
end if;
if first_state_sram_input_id = 11219 then
	sram_write <= x"D0626000";
end if;
if first_state_sram_input_id = 11220 then
	sram_write <= x"C0660000";
end if;
if first_state_sram_input_id = 11221 then
	sram_write <= x"44202000";
end if;
if first_state_sram_input_id = 11222 then
	sram_write <= x"CCA60000";
end if;
if first_state_sram_input_id = 11223 then
	sram_write <= x"CC860004";
end if;
if first_state_sram_input_id = 11224 then
	sram_write <= x"CC260008";
end if;
if first_state_sram_input_id = 11225 then
	sram_write <= x"02640029";
end if;
if first_state_sram_input_id = 11226 then
	sram_write <= x"22660220";
end if;
if first_state_sram_input_id = 11227 then
	sram_write <= x"D0626000";
end if;
if first_state_sram_input_id = 11228 then
	sram_write <= x"C0660000";
end if;
if first_state_sram_input_id = 11229 then
	sram_write <= x"CCA60000";
end if;
if first_state_sram_input_id = 11230 then
	sram_write <= x"CC260004";
end if;
if first_state_sram_input_id = 11231 then
	sram_write <= x"CC660008";
end if;
if first_state_sram_input_id = 11232 then
	sram_write <= x"02440051";
end if;
if first_state_sram_input_id = 11233 then
	sram_write <= x"22440220";
end if;
if first_state_sram_input_id = 11234 then
	sram_write <= x"D0224000";
end if;
if first_state_sram_input_id = 11235 then
	sram_write <= x"C0220000";
end if;
if first_state_sram_input_id = 11236 then
	sram_write <= x"CC220000";
end if;
if first_state_sram_input_id = 11237 then
	sram_write <= x"CC420004";
end if;
if first_state_sram_input_id = 11238 then
	sram_write <= x"CC620008";
end if;
if first_state_sram_input_id = 11239 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 11240 then
	sram_write <= x"48244000";
end if;
if first_state_sram_input_id = 11241 then
	sram_write <= x"C840001C";
end if;
if first_state_sram_input_id = 11242 then
	sram_write <= x"40224000";
end if;
if first_state_sram_input_id = 11243 then
	sram_write <= x"C47C0000";
end if;
if first_state_sram_input_id = 11244 then
	sram_write <= x"C45C0004";
end if;
if first_state_sram_input_id = 11245 then
	sram_write <= x"CC9C0030";
end if;
if first_state_sram_input_id = 11246 then
	sram_write <= x"CC5C0038";
end if;
if first_state_sram_input_id = 11247 then
	sram_write <= x"C43C0040";
end if;
if first_state_sram_input_id = 11248 then
	sram_write <= x"CC7C0048";
end if;
if first_state_sram_input_id = 11249 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11250 then
	sram_write <= x"03DC0058";
end if;
if first_state_sram_input_id = 11251 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11252 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11253 then
	sram_write <= x"8200083C";
end if;
if first_state_sram_input_id = 11254 then
	sram_write <= x"07DC0058";
end if;
if first_state_sram_input_id = 11255 then
	sram_write <= x"CC3C0050";
end if;
if first_state_sram_input_id = 11256 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11257 then
	sram_write <= x"03DC0060";
end if;
if first_state_sram_input_id = 11258 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11259 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11260 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 11261 then
	sram_write <= x"07DC0060";
end if;
if first_state_sram_input_id = 11262 then
	sram_write <= x"C8400068";
end if;
if first_state_sram_input_id = 11263 then
	sram_write <= x"48642000";
end if;
if first_state_sram_input_id = 11264 then
	sram_write <= x"C8800064";
end if;
if first_state_sram_input_id = 11265 then
	sram_write <= x"44668000";
end if;
if first_state_sram_input_id = 11266 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 11267 then
	sram_write <= x"C8A00060";
end if;
if first_state_sram_input_id = 11268 then
	sram_write <= x"4466A000";
end if;
if first_state_sram_input_id = 11269 then
	sram_write <= x"48662000";
end if;
if first_state_sram_input_id = 11270 then
	sram_write <= x"C8C0005C";
end if;
if first_state_sram_input_id = 11271 then
	sram_write <= x"4066C000";
end if;
if first_state_sram_input_id = 11272 then
	sram_write <= x"48262000";
end if;
if first_state_sram_input_id = 11273 then
	sram_write <= x"C8600058";
end if;
if first_state_sram_input_id = 11274 then
	sram_write <= x"44226000";
end if;
if first_state_sram_input_id = 11275 then
	sram_write <= x"C8FC0048";
end if;
if first_state_sram_input_id = 11276 then
	sram_write <= x"4822E000";
end if;
if first_state_sram_input_id = 11277 then
	sram_write <= x"C9000098";
end if;
if first_state_sram_input_id = 11278 then
	sram_write <= x"CC7C0058";
end if;
if first_state_sram_input_id = 11279 then
	sram_write <= x"CCDC0060";
end if;
if first_state_sram_input_id = 11280 then
	sram_write <= x"CCBC0068";
end if;
if first_state_sram_input_id = 11281 then
	sram_write <= x"CC9C0070";
end if;
if first_state_sram_input_id = 11282 then
	sram_write <= x"CC5C0078";
end if;
if first_state_sram_input_id = 11283 then
	sram_write <= x"CD1C0080";
end if;
if first_state_sram_input_id = 11284 then
	sram_write <= x"CC3C0088";
end if;
if first_state_sram_input_id = 11285 then
	sram_write <= x"8E30B07C";
end if;
if first_state_sram_input_id = 11286 then
	sram_write <= x"45230000";
end if;
if first_state_sram_input_id = 11287 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11288 then
	sram_write <= x"40212000";
end if;
if first_state_sram_input_id = 11289 then
	sram_write <= x"03DC0098";
end if;
if first_state_sram_input_id = 11290 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11291 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11292 then
	sram_write <= x"82000EC4";
end if;
if first_state_sram_input_id = 11293 then
	sram_write <= x"07DC0098";
end if;
if first_state_sram_input_id = 11294 then
	sram_write <= x"8200B0E8";
end if;
if first_state_sram_input_id = 11295 then
	sram_write <= x"8E02B0CC";
end if;
if first_state_sram_input_id = 11296 then
	sram_write <= x"C9200090";
end if;
if first_state_sram_input_id = 11297 then
	sram_write <= x"8F22B0AC";
end if;
if first_state_sram_input_id = 11298 then
	sram_write <= x"41230000";
end if;
if first_state_sram_input_id = 11299 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11300 then
	sram_write <= x"40212000";
end if;
if first_state_sram_input_id = 11301 then
	sram_write <= x"03DC0098";
end if;
if first_state_sram_input_id = 11302 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11303 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11304 then
	sram_write <= x"82000EC4";
end if;
if first_state_sram_input_id = 11305 then
	sram_write <= x"07DC0098";
end if;
if first_state_sram_input_id = 11306 then
	sram_write <= x"8200B0C8";
end if;
if first_state_sram_input_id = 11307 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 11308 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11309 then
	sram_write <= x"03DC0098";
end if;
if first_state_sram_input_id = 11310 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11311 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11312 then
	sram_write <= x"8200084C";
end if;
if first_state_sram_input_id = 11313 then
	sram_write <= x"07DC0098";
end if;
if first_state_sram_input_id = 11314 then
	sram_write <= x"8200B0E8";
end if;
if first_state_sram_input_id = 11315 then
	sram_write <= x"0220FFFF";
end if;
if first_state_sram_input_id = 11316 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11317 then
	sram_write <= x"03DC0098";
end if;
if first_state_sram_input_id = 11318 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11319 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11320 then
	sram_write <= x"8200084C";
end if;
if first_state_sram_input_id = 11321 then
	sram_write <= x"07DC0098";
end if;
if first_state_sram_input_id = 11322 then
	sram_write <= x"C85C0080";
end if;
if first_state_sram_input_id = 11323 then
	sram_write <= x"C87C0088";
end if;
if first_state_sram_input_id = 11324 then
	sram_write <= x"CC3C0090";
end if;
if first_state_sram_input_id = 11325 then
	sram_write <= x"8E64B11C";
end if;
if first_state_sram_input_id = 11326 then
	sram_write <= x"44664000";
end if;
if first_state_sram_input_id = 11327 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11328 then
	sram_write <= x"40206000";
end if;
if first_state_sram_input_id = 11329 then
	sram_write <= x"03DC00A0";
end if;
if first_state_sram_input_id = 11330 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11331 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11332 then
	sram_write <= x"82001270";
end if;
if first_state_sram_input_id = 11333 then
	sram_write <= x"07DC00A0";
end if;
if first_state_sram_input_id = 11334 then
	sram_write <= x"8200B190";
end if;
if first_state_sram_input_id = 11335 then
	sram_write <= x"8E06B170";
end if;
if first_state_sram_input_id = 11336 then
	sram_write <= x"C8800090";
end if;
if first_state_sram_input_id = 11337 then
	sram_write <= x"8E86B14C";
end if;
if first_state_sram_input_id = 11338 then
	sram_write <= x"40664000";
end if;
if first_state_sram_input_id = 11339 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11340 then
	sram_write <= x"40206000";
end if;
if first_state_sram_input_id = 11341 then
	sram_write <= x"03DC00A0";
end if;
if first_state_sram_input_id = 11342 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11343 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11344 then
	sram_write <= x"82001270";
end if;
if first_state_sram_input_id = 11345 then
	sram_write <= x"07DC00A0";
end if;
if first_state_sram_input_id = 11346 then
	sram_write <= x"8200B16C";
end if;
if first_state_sram_input_id = 11347 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 11348 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11349 then
	sram_write <= x"40206000";
end if;
if first_state_sram_input_id = 11350 then
	sram_write <= x"03DC00A0";
end if;
if first_state_sram_input_id = 11351 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11352 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11353 then
	sram_write <= x"82000B88";
end if;
if first_state_sram_input_id = 11354 then
	sram_write <= x"07DC00A0";
end if;
if first_state_sram_input_id = 11355 then
	sram_write <= x"8200B190";
end if;
if first_state_sram_input_id = 11356 then
	sram_write <= x"0220FFFF";
end if;
if first_state_sram_input_id = 11357 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11358 then
	sram_write <= x"40206000";
end if;
if first_state_sram_input_id = 11359 then
	sram_write <= x"03DC00A0";
end if;
if first_state_sram_input_id = 11360 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11361 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11362 then
	sram_write <= x"82000B88";
end if;
if first_state_sram_input_id = 11363 then
	sram_write <= x"07DC00A0";
end if;
if first_state_sram_input_id = 11364 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11365 then
	sram_write <= x"03DC00A0";
end if;
if first_state_sram_input_id = 11366 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11367 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11368 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 11369 then
	sram_write <= x"07DC00A0";
end if;
if first_state_sram_input_id = 11370 then
	sram_write <= x"C85C0090";
end if;
if first_state_sram_input_id = 11371 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 11372 then
	sram_write <= x"C85C0050";
end if;
if first_state_sram_input_id = 11373 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 11374 then
	sram_write <= x"C03C0040";
end if;
if first_state_sram_input_id = 11375 then
	sram_write <= x"02220001";
end if;
if first_state_sram_input_id = 11376 then
	sram_write <= x"48422000";
end if;
if first_state_sram_input_id = 11377 then
	sram_write <= x"C87C0038";
end if;
if first_state_sram_input_id = 11378 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 11379 then
	sram_write <= x"CC3C0098";
end if;
if first_state_sram_input_id = 11380 then
	sram_write <= x"C43C00A0";
end if;
if first_state_sram_input_id = 11381 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11382 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 11383 then
	sram_write <= x"03DC00AC";
end if;
if first_state_sram_input_id = 11384 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11385 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11386 then
	sram_write <= x"8200083C";
end if;
if first_state_sram_input_id = 11387 then
	sram_write <= x"07DC00AC";
end if;
if first_state_sram_input_id = 11388 then
	sram_write <= x"CC3C00A8";
end if;
if first_state_sram_input_id = 11389 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11390 then
	sram_write <= x"03DC00B8";
end if;
if first_state_sram_input_id = 11391 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11392 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11393 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 11394 then
	sram_write <= x"07DC00B8";
end if;
if first_state_sram_input_id = 11395 then
	sram_write <= x"C85C0078";
end if;
if first_state_sram_input_id = 11396 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 11397 then
	sram_write <= x"C87C0070";
end if;
if first_state_sram_input_id = 11398 then
	sram_write <= x"44446000";
end if;
if first_state_sram_input_id = 11399 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 11400 then
	sram_write <= x"C87C0068";
end if;
if first_state_sram_input_id = 11401 then
	sram_write <= x"44446000";
end if;
if first_state_sram_input_id = 11402 then
	sram_write <= x"48442000";
end if;
if first_state_sram_input_id = 11403 then
	sram_write <= x"C87C0060";
end if;
if first_state_sram_input_id = 11404 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 11405 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 11406 then
	sram_write <= x"C85C0058";
end if;
if first_state_sram_input_id = 11407 then
	sram_write <= x"44224000";
end if;
if first_state_sram_input_id = 11408 then
	sram_write <= x"C85C0030";
end if;
if first_state_sram_input_id = 11409 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 11410 then
	sram_write <= x"C87C0080";
end if;
if first_state_sram_input_id = 11411 then
	sram_write <= x"CC3C00B0";
end if;
if first_state_sram_input_id = 11412 then
	sram_write <= x"8E26B278";
end if;
if first_state_sram_input_id = 11413 then
	sram_write <= x"44826000";
end if;
if first_state_sram_input_id = 11414 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11415 then
	sram_write <= x"40208000";
end if;
if first_state_sram_input_id = 11416 then
	sram_write <= x"03DC00C0";
end if;
if first_state_sram_input_id = 11417 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11418 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11419 then
	sram_write <= x"82000EC4";
end if;
if first_state_sram_input_id = 11420 then
	sram_write <= x"07DC00C0";
end if;
if first_state_sram_input_id = 11421 then
	sram_write <= x"8200B2E4";
end if;
if first_state_sram_input_id = 11422 then
	sram_write <= x"8E02B2C8";
end if;
if first_state_sram_input_id = 11423 then
	sram_write <= x"C8800090";
end if;
if first_state_sram_input_id = 11424 then
	sram_write <= x"8E82B2A8";
end if;
if first_state_sram_input_id = 11425 then
	sram_write <= x"40826000";
end if;
if first_state_sram_input_id = 11426 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11427 then
	sram_write <= x"40208000";
end if;
if first_state_sram_input_id = 11428 then
	sram_write <= x"03DC00C0";
end if;
if first_state_sram_input_id = 11429 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11430 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11431 then
	sram_write <= x"82000EC4";
end if;
if first_state_sram_input_id = 11432 then
	sram_write <= x"07DC00C0";
end if;
if first_state_sram_input_id = 11433 then
	sram_write <= x"8200B2C4";
end if;
if first_state_sram_input_id = 11434 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 11435 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11436 then
	sram_write <= x"03DC00C0";
end if;
if first_state_sram_input_id = 11437 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11438 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11439 then
	sram_write <= x"8200084C";
end if;
if first_state_sram_input_id = 11440 then
	sram_write <= x"07DC00C0";
end if;
if first_state_sram_input_id = 11441 then
	sram_write <= x"8200B2E4";
end if;
if first_state_sram_input_id = 11442 then
	sram_write <= x"0220FFFF";
end if;
if first_state_sram_input_id = 11443 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11444 then
	sram_write <= x"03DC00C0";
end if;
if first_state_sram_input_id = 11445 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11446 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11447 then
	sram_write <= x"8200084C";
end if;
if first_state_sram_input_id = 11448 then
	sram_write <= x"07DC00C0";
end if;
if first_state_sram_input_id = 11449 then
	sram_write <= x"C85C0080";
end if;
if first_state_sram_input_id = 11450 then
	sram_write <= x"C87C00B0";
end if;
if first_state_sram_input_id = 11451 then
	sram_write <= x"CC3C00B8";
end if;
if first_state_sram_input_id = 11452 then
	sram_write <= x"8E64B318";
end if;
if first_state_sram_input_id = 11453 then
	sram_write <= x"44464000";
end if;
if first_state_sram_input_id = 11454 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11455 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 11456 then
	sram_write <= x"03DC00C8";
end if;
if first_state_sram_input_id = 11457 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11458 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11459 then
	sram_write <= x"82001270";
end if;
if first_state_sram_input_id = 11460 then
	sram_write <= x"07DC00C8";
end if;
if first_state_sram_input_id = 11461 then
	sram_write <= x"8200B38C";
end if;
if first_state_sram_input_id = 11462 then
	sram_write <= x"8E06B36C";
end if;
if first_state_sram_input_id = 11463 then
	sram_write <= x"C8800090";
end if;
if first_state_sram_input_id = 11464 then
	sram_write <= x"8E86B348";
end if;
if first_state_sram_input_id = 11465 then
	sram_write <= x"40464000";
end if;
if first_state_sram_input_id = 11466 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11467 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 11468 then
	sram_write <= x"03DC00C8";
end if;
if first_state_sram_input_id = 11469 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11470 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11471 then
	sram_write <= x"82001270";
end if;
if first_state_sram_input_id = 11472 then
	sram_write <= x"07DC00C8";
end if;
if first_state_sram_input_id = 11473 then
	sram_write <= x"8200B368";
end if;
if first_state_sram_input_id = 11474 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 11475 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11476 then
	sram_write <= x"40206000";
end if;
if first_state_sram_input_id = 11477 then
	sram_write <= x"03DC00C8";
end if;
if first_state_sram_input_id = 11478 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11479 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11480 then
	sram_write <= x"82000B88";
end if;
if first_state_sram_input_id = 11481 then
	sram_write <= x"07DC00C8";
end if;
if first_state_sram_input_id = 11482 then
	sram_write <= x"8200B38C";
end if;
if first_state_sram_input_id = 11483 then
	sram_write <= x"0220FFFF";
end if;
if first_state_sram_input_id = 11484 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11485 then
	sram_write <= x"40206000";
end if;
if first_state_sram_input_id = 11486 then
	sram_write <= x"03DC00C8";
end if;
if first_state_sram_input_id = 11487 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11488 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11489 then
	sram_write <= x"82000B88";
end if;
if first_state_sram_input_id = 11490 then
	sram_write <= x"07DC00C8";
end if;
if first_state_sram_input_id = 11491 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11492 then
	sram_write <= x"03DC00C8";
end if;
if first_state_sram_input_id = 11493 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11494 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11495 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 11496 then
	sram_write <= x"07DC00C8";
end if;
if first_state_sram_input_id = 11497 then
	sram_write <= x"C85C00B8";
end if;
if first_state_sram_input_id = 11498 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 11499 then
	sram_write <= x"C85C00A8";
end if;
if first_state_sram_input_id = 11500 then
	sram_write <= x"48424000";
end if;
if first_state_sram_input_id = 11501 then
	sram_write <= x"C83C0098";
end if;
if first_state_sram_input_id = 11502 then
	sram_write <= x"C87C0048";
end if;
if first_state_sram_input_id = 11503 then
	sram_write <= x"C89C0030";
end if;
if first_state_sram_input_id = 11504 then
	sram_write <= x"C03C00A0";
end if;
if first_state_sram_input_id = 11505 then
	sram_write <= x"C05C0004";
end if;
if first_state_sram_input_id = 11506 then
	sram_write <= x"C07C0000";
end if;
if first_state_sram_input_id = 11507 then
	sram_write <= x"8200AE14";
end if;
if first_state_sram_input_id = 11508 then
	sram_write <= x"8620B570";
end if;
if first_state_sram_input_id = 11509 then
	sram_write <= x"58420000";
end if;
if first_state_sram_input_id = 11510 then
	sram_write <= x"C8600010";
end if;
if first_state_sram_input_id = 11511 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 11512 then
	sram_write <= x"C880000C";
end if;
if first_state_sram_input_id = 11513 then
	sram_write <= x"44A48000";
end if;
if first_state_sram_input_id = 11514 then
	sram_write <= x"02800000";
end if;
if first_state_sram_input_id = 11515 then
	sram_write <= x"40C00000";
end if;
if first_state_sram_input_id = 11516 then
	sram_write <= x"CC9C0000";
end if;
if first_state_sram_input_id = 11517 then
	sram_write <= x"CC7C0008";
end if;
if first_state_sram_input_id = 11518 then
	sram_write <= x"C43C0010";
end if;
if first_state_sram_input_id = 11519 then
	sram_write <= x"CC3C0018";
end if;
if first_state_sram_input_id = 11520 then
	sram_write <= x"CCDC0020";
end if;
if first_state_sram_input_id = 11521 then
	sram_write <= x"C45C0028";
end if;
if first_state_sram_input_id = 11522 then
	sram_write <= x"C47C002C";
end if;
if first_state_sram_input_id = 11523 then
	sram_write <= x"CC5C0030";
end if;
if first_state_sram_input_id = 11524 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11525 then
	sram_write <= x"00280000";
end if;
if first_state_sram_input_id = 11526 then
	sram_write <= x"40802000";
end if;
if first_state_sram_input_id = 11527 then
	sram_write <= x"4060A000";
end if;
if first_state_sram_input_id = 11528 then
	sram_write <= x"4040C000";
end if;
if first_state_sram_input_id = 11529 then
	sram_write <= x"4020C000";
end if;
if first_state_sram_input_id = 11530 then
	sram_write <= x"03DC0040";
end if;
if first_state_sram_input_id = 11531 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11532 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11533 then
	sram_write <= x"8200AE14";
end if;
if first_state_sram_input_id = 11534 then
	sram_write <= x"07DC0040";
end if;
if first_state_sram_input_id = 11535 then
	sram_write <= x"C820001C";
end if;
if first_state_sram_input_id = 11536 then
	sram_write <= x"C85C0030";
end if;
if first_state_sram_input_id = 11537 then
	sram_write <= x"40642000";
end if;
if first_state_sram_input_id = 11538 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 11539 then
	sram_write <= x"C05C002C";
end if;
if first_state_sram_input_id = 11540 then
	sram_write <= x"02640002";
end if;
if first_state_sram_input_id = 11541 then
	sram_write <= x"C85C0020";
end if;
if first_state_sram_input_id = 11542 then
	sram_write <= x"C89C0018";
end if;
if first_state_sram_input_id = 11543 then
	sram_write <= x"C09C0028";
end if;
if first_state_sram_input_id = 11544 then
	sram_write <= x"CC3C0038";
end if;
if first_state_sram_input_id = 11545 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11546 then
	sram_write <= x"00480000";
end if;
if first_state_sram_input_id = 11547 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 11548 then
	sram_write <= x"03DC0048";
end if;
if first_state_sram_input_id = 11549 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11550 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11551 then
	sram_write <= x"8200AE14";
end if;
if first_state_sram_input_id = 11552 then
	sram_write <= x"07DC0048";
end if;
if first_state_sram_input_id = 11553 then
	sram_write <= x"C03C0010";
end if;
if first_state_sram_input_id = 11554 then
	sram_write <= x"06220001";
end if;
if first_state_sram_input_id = 11555 then
	sram_write <= x"C05C0028";
end if;
if first_state_sram_input_id = 11556 then
	sram_write <= x"02440001";
end if;
if first_state_sram_input_id = 11557 then
	sram_write <= x"02600005";
end if;
if first_state_sram_input_id = 11558 then
	sram_write <= x"8646B4A4";
end if;
if first_state_sram_input_id = 11559 then
	sram_write <= x"06440005";
end if;
if first_state_sram_input_id = 11560 then
	sram_write <= x"8200B4A4";
end if;
if first_state_sram_input_id = 11561 then
	sram_write <= x"8620B56C";
end if;
if first_state_sram_input_id = 11562 then
	sram_write <= x"58220000";
end if;
if first_state_sram_input_id = 11563 then
	sram_write <= x"C85C0008";
end if;
if first_state_sram_input_id = 11564 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 11565 then
	sram_write <= x"C85C0000";
end if;
if first_state_sram_input_id = 11566 then
	sram_write <= x"44624000";
end if;
if first_state_sram_input_id = 11567 then
	sram_write <= x"02600000";
end if;
if first_state_sram_input_id = 11568 then
	sram_write <= x"C85C0020";
end if;
if first_state_sram_input_id = 11569 then
	sram_write <= x"C89C0018";
end if;
if first_state_sram_input_id = 11570 then
	sram_write <= x"C09C002C";
end if;
if first_state_sram_input_id = 11571 then
	sram_write <= x"C43C0040";
end if;
if first_state_sram_input_id = 11572 then
	sram_write <= x"C45C0044";
end if;
if first_state_sram_input_id = 11573 then
	sram_write <= x"CC3C0048";
end if;
if first_state_sram_input_id = 11574 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11575 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 11576 then
	sram_write <= x"00680000";
end if;
if first_state_sram_input_id = 11577 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 11578 then
	sram_write <= x"03DC0058";
end if;
if first_state_sram_input_id = 11579 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11580 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11581 then
	sram_write <= x"8200AE14";
end if;
if first_state_sram_input_id = 11582 then
	sram_write <= x"07DC0058";
end if;
if first_state_sram_input_id = 11583 then
	sram_write <= x"C83C0038";
end if;
if first_state_sram_input_id = 11584 then
	sram_write <= x"C85C0048";
end if;
if first_state_sram_input_id = 11585 then
	sram_write <= x"40642000";
end if;
if first_state_sram_input_id = 11586 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 11587 then
	sram_write <= x"C05C002C";
end if;
if first_state_sram_input_id = 11588 then
	sram_write <= x"02640002";
end if;
if first_state_sram_input_id = 11589 then
	sram_write <= x"C83C0020";
end if;
if first_state_sram_input_id = 11590 then
	sram_write <= x"C89C0018";
end if;
if first_state_sram_input_id = 11591 then
	sram_write <= x"C09C0044";
end if;
if first_state_sram_input_id = 11592 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11593 then
	sram_write <= x"00480000";
end if;
if first_state_sram_input_id = 11594 then
	sram_write <= x"40402000";
end if;
if first_state_sram_input_id = 11595 then
	sram_write <= x"03DC0058";
end if;
if first_state_sram_input_id = 11596 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11597 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11598 then
	sram_write <= x"8200AE14";
end if;
if first_state_sram_input_id = 11599 then
	sram_write <= x"07DC0058";
end if;
if first_state_sram_input_id = 11600 then
	sram_write <= x"C03C0040";
end if;
if first_state_sram_input_id = 11601 then
	sram_write <= x"06220001";
end if;
if first_state_sram_input_id = 11602 then
	sram_write <= x"C05C0044";
end if;
if first_state_sram_input_id = 11603 then
	sram_write <= x"02440001";
end if;
if first_state_sram_input_id = 11604 then
	sram_write <= x"02600005";
end if;
if first_state_sram_input_id = 11605 then
	sram_write <= x"8646B560";
end if;
if first_state_sram_input_id = 11606 then
	sram_write <= x"06440005";
end if;
if first_state_sram_input_id = 11607 then
	sram_write <= x"8200B560";
end if;
if first_state_sram_input_id = 11608 then
	sram_write <= x"C83C0018";
end if;
if first_state_sram_input_id = 11609 then
	sram_write <= x"C07C002C";
end if;
if first_state_sram_input_id = 11610 then
	sram_write <= x"8200B3D0";
end if;
if first_state_sram_input_id = 11611 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 11612 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 11613 then
	sram_write <= x"8620B6F8";
end if;
if first_state_sram_input_id = 11614 then
	sram_write <= x"58220000";
end if;
if first_state_sram_input_id = 11615 then
	sram_write <= x"C8400010";
end if;
if first_state_sram_input_id = 11616 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 11617 then
	sram_write <= x"C860000C";
end if;
if first_state_sram_input_id = 11618 then
	sram_write <= x"44826000";
end if;
if first_state_sram_input_id = 11619 then
	sram_write <= x"C8200008";
end if;
if first_state_sram_input_id = 11620 then
	sram_write <= x"02800000";
end if;
if first_state_sram_input_id = 11621 then
	sram_write <= x"40A00000";
end if;
if first_state_sram_input_id = 11622 then
	sram_write <= x"CC5C0000";
end if;
if first_state_sram_input_id = 11623 then
	sram_write <= x"C43C0008";
end if;
if first_state_sram_input_id = 11624 then
	sram_write <= x"CC9C0010";
end if;
if first_state_sram_input_id = 11625 then
	sram_write <= x"CC7C0018";
end if;
if first_state_sram_input_id = 11626 then
	sram_write <= x"CCBC0020";
end if;
if first_state_sram_input_id = 11627 then
	sram_write <= x"C45C0028";
end if;
if first_state_sram_input_id = 11628 then
	sram_write <= x"C47C002C";
end if;
if first_state_sram_input_id = 11629 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11630 then
	sram_write <= x"00280000";
end if;
if first_state_sram_input_id = 11631 then
	sram_write <= x"40602000";
end if;
if first_state_sram_input_id = 11632 then
	sram_write <= x"4040A000";
end if;
if first_state_sram_input_id = 11633 then
	sram_write <= x"4020A000";
end if;
if first_state_sram_input_id = 11634 then
	sram_write <= x"03DC0038";
end if;
if first_state_sram_input_id = 11635 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11636 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11637 then
	sram_write <= x"8200AE14";
end if;
if first_state_sram_input_id = 11638 then
	sram_write <= x"07DC0038";
end if;
if first_state_sram_input_id = 11639 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 11640 then
	sram_write <= x"C05C002C";
end if;
if first_state_sram_input_id = 11641 then
	sram_write <= x"02640002";
end if;
if first_state_sram_input_id = 11642 then
	sram_write <= x"C83C0020";
end if;
if first_state_sram_input_id = 11643 then
	sram_write <= x"C87C0018";
end if;
if first_state_sram_input_id = 11644 then
	sram_write <= x"C89C0010";
end if;
if first_state_sram_input_id = 11645 then
	sram_write <= x"C09C0028";
end if;
if first_state_sram_input_id = 11646 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11647 then
	sram_write <= x"00480000";
end if;
if first_state_sram_input_id = 11648 then
	sram_write <= x"40402000";
end if;
if first_state_sram_input_id = 11649 then
	sram_write <= x"03DC0038";
end if;
if first_state_sram_input_id = 11650 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11651 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11652 then
	sram_write <= x"8200AE14";
end if;
if first_state_sram_input_id = 11653 then
	sram_write <= x"07DC0038";
end if;
if first_state_sram_input_id = 11654 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 11655 then
	sram_write <= x"C05C0028";
end if;
if first_state_sram_input_id = 11656 then
	sram_write <= x"02640001";
end if;
if first_state_sram_input_id = 11657 then
	sram_write <= x"02800005";
end if;
if first_state_sram_input_id = 11658 then
	sram_write <= x"8668B634";
end if;
if first_state_sram_input_id = 11659 then
	sram_write <= x"06660005";
end if;
if first_state_sram_input_id = 11660 then
	sram_write <= x"8200B634";
end if;
if first_state_sram_input_id = 11661 then
	sram_write <= x"C83C0010";
end if;
if first_state_sram_input_id = 11662 then
	sram_write <= x"C09C002C";
end if;
if first_state_sram_input_id = 11663 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11664 then
	sram_write <= x"00460000";
end if;
if first_state_sram_input_id = 11665 then
	sram_write <= x"00680000";
end if;
if first_state_sram_input_id = 11666 then
	sram_write <= x"03DC0038";
end if;
if first_state_sram_input_id = 11667 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11668 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11669 then
	sram_write <= x"8200B3D0";
end if;
if first_state_sram_input_id = 11670 then
	sram_write <= x"07DC0038";
end if;
if first_state_sram_input_id = 11671 then
	sram_write <= x"C03C0008";
end if;
if first_state_sram_input_id = 11672 then
	sram_write <= x"06220001";
end if;
if first_state_sram_input_id = 11673 then
	sram_write <= x"C05C0028";
end if;
if first_state_sram_input_id = 11674 then
	sram_write <= x"02440002";
end if;
if first_state_sram_input_id = 11675 then
	sram_write <= x"02600005";
end if;
if first_state_sram_input_id = 11676 then
	sram_write <= x"8646B67C";
end if;
if first_state_sram_input_id = 11677 then
	sram_write <= x"06440005";
end if;
if first_state_sram_input_id = 11678 then
	sram_write <= x"8200B67C";
end if;
if first_state_sram_input_id = 11679 then
	sram_write <= x"C07C002C";
end if;
if first_state_sram_input_id = 11680 then
	sram_write <= x"02660004";
end if;
if first_state_sram_input_id = 11681 then
	sram_write <= x"8620B6F4";
end if;
if first_state_sram_input_id = 11682 then
	sram_write <= x"58220000";
end if;
if first_state_sram_input_id = 11683 then
	sram_write <= x"C85C0000";
end if;
if first_state_sram_input_id = 11684 then
	sram_write <= x"48224000";
end if;
if first_state_sram_input_id = 11685 then
	sram_write <= x"C85C0018";
end if;
if first_state_sram_input_id = 11686 then
	sram_write <= x"44224000";
end if;
if first_state_sram_input_id = 11687 then
	sram_write <= x"02800004";
end if;
if first_state_sram_input_id = 11688 then
	sram_write <= x"C47C0030";
end if;
if first_state_sram_input_id = 11689 then
	sram_write <= x"C45C0034";
end if;
if first_state_sram_input_id = 11690 then
	sram_write <= x"C43C0038";
end if;
if first_state_sram_input_id = 11691 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11692 then
	sram_write <= x"00280000";
end if;
if first_state_sram_input_id = 11693 then
	sram_write <= x"03DC0044";
end if;
if first_state_sram_input_id = 11694 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11695 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11696 then
	sram_write <= x"8200B3D0";
end if;
if first_state_sram_input_id = 11697 then
	sram_write <= x"07DC0044";
end if;
if first_state_sram_input_id = 11698 then
	sram_write <= x"C03C0038";
end if;
if first_state_sram_input_id = 11699 then
	sram_write <= x"06220001";
end if;
if first_state_sram_input_id = 11700 then
	sram_write <= x"C05C0034";
end if;
if first_state_sram_input_id = 11701 then
	sram_write <= x"02440002";
end if;
if first_state_sram_input_id = 11702 then
	sram_write <= x"02600005";
end if;
if first_state_sram_input_id = 11703 then
	sram_write <= x"8646B6E8";
end if;
if first_state_sram_input_id = 11704 then
	sram_write <= x"06440005";
end if;
if first_state_sram_input_id = 11705 then
	sram_write <= x"8200B6E8";
end if;
if first_state_sram_input_id = 11706 then
	sram_write <= x"C07C0030";
end if;
if first_state_sram_input_id = 11707 then
	sram_write <= x"02660004";
end if;
if first_state_sram_input_id = 11708 then
	sram_write <= x"8200B574";
end if;
if first_state_sram_input_id = 11709 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 11710 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 11711 then
	sram_write <= x"8640B928";
end if;
if first_state_sram_input_id = 11712 then
	sram_write <= x"02600003";
end if;
if first_state_sram_input_id = 11713 then
	sram_write <= x"40200000";
end if;
if first_state_sram_input_id = 11714 then
	sram_write <= x"CC3C0000";
end if;
if first_state_sram_input_id = 11715 then
	sram_write <= x"C43C0008";
end if;
if first_state_sram_input_id = 11716 then
	sram_write <= x"C45C000C";
end if;
if first_state_sram_input_id = 11717 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11718 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 11719 then
	sram_write <= x"03DC0018";
end if;
if first_state_sram_input_id = 11720 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11721 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11722 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 11723 then
	sram_write <= x"07DC0018";
end if;
if first_state_sram_input_id = 11724 then
	sram_write <= x"00420000";
end if;
if first_state_sram_input_id = 11725 then
	sram_write <= x"022000C4";
end if;
if first_state_sram_input_id = 11726 then
	sram_write <= x"C0620000";
end if;
if first_state_sram_input_id = 11727 then
	sram_write <= x"C43C0010";
end if;
if first_state_sram_input_id = 11728 then
	sram_write <= x"C45C0014";
end if;
if first_state_sram_input_id = 11729 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11730 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 11731 then
	sram_write <= x"03DC0020";
end if;
if first_state_sram_input_id = 11732 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11733 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11734 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 11735 then
	sram_write <= x"07DC0020";
end if;
if first_state_sram_input_id = 11736 then
	sram_write <= x"005A0000";
end if;
if first_state_sram_input_id = 11737 then
	sram_write <= x"03BA0008";
end if;
if first_state_sram_input_id = 11738 then
	sram_write <= x"C4240004";
end if;
if first_state_sram_input_id = 11739 then
	sram_write <= x"C03C0014";
end if;
if first_state_sram_input_id = 11740 then
	sram_write <= x"C4240000";
end if;
if first_state_sram_input_id = 11741 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 11742 then
	sram_write <= x"C05C000C";
end if;
if first_state_sram_input_id = 11743 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 11744 then
	sram_write <= x"C09C0008";
end if;
if first_state_sram_input_id = 11745 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 11746 then
	sram_write <= x"06240001";
end if;
if first_state_sram_input_id = 11747 then
	sram_write <= x"8620B924";
end if;
if first_state_sram_input_id = 11748 then
	sram_write <= x"02400003";
end if;
if first_state_sram_input_id = 11749 then
	sram_write <= x"C83C0000";
end if;
if first_state_sram_input_id = 11750 then
	sram_write <= x"C43C0018";
end if;
if first_state_sram_input_id = 11751 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11752 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 11753 then
	sram_write <= x"03DC0024";
end if;
if first_state_sram_input_id = 11754 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11755 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11756 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 11757 then
	sram_write <= x"07DC0024";
end if;
if first_state_sram_input_id = 11758 then
	sram_write <= x"00420000";
end if;
if first_state_sram_input_id = 11759 then
	sram_write <= x"C03C0010";
end if;
if first_state_sram_input_id = 11760 then
	sram_write <= x"C0620000";
end if;
if first_state_sram_input_id = 11761 then
	sram_write <= x"C45C001C";
end if;
if first_state_sram_input_id = 11762 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11763 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 11764 then
	sram_write <= x"03DC0028";
end if;
if first_state_sram_input_id = 11765 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11766 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11767 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 11768 then
	sram_write <= x"07DC0028";
end if;
if first_state_sram_input_id = 11769 then
	sram_write <= x"005A0000";
end if;
if first_state_sram_input_id = 11770 then
	sram_write <= x"03BA0008";
end if;
if first_state_sram_input_id = 11771 then
	sram_write <= x"C4240004";
end if;
if first_state_sram_input_id = 11772 then
	sram_write <= x"C03C001C";
end if;
if first_state_sram_input_id = 11773 then
	sram_write <= x"C4240000";
end if;
if first_state_sram_input_id = 11774 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 11775 then
	sram_write <= x"C05C0018";
end if;
if first_state_sram_input_id = 11776 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 11777 then
	sram_write <= x"C09C0008";
end if;
if first_state_sram_input_id = 11778 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 11779 then
	sram_write <= x"06240001";
end if;
if first_state_sram_input_id = 11780 then
	sram_write <= x"8620B920";
end if;
if first_state_sram_input_id = 11781 then
	sram_write <= x"02400003";
end if;
if first_state_sram_input_id = 11782 then
	sram_write <= x"C83C0000";
end if;
if first_state_sram_input_id = 11783 then
	sram_write <= x"C43C0020";
end if;
if first_state_sram_input_id = 11784 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11785 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 11786 then
	sram_write <= x"03DC002C";
end if;
if first_state_sram_input_id = 11787 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11788 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11789 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 11790 then
	sram_write <= x"07DC002C";
end if;
if first_state_sram_input_id = 11791 then
	sram_write <= x"00420000";
end if;
if first_state_sram_input_id = 11792 then
	sram_write <= x"C03C0010";
end if;
if first_state_sram_input_id = 11793 then
	sram_write <= x"C0620000";
end if;
if first_state_sram_input_id = 11794 then
	sram_write <= x"C45C0024";
end if;
if first_state_sram_input_id = 11795 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11796 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 11797 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 11798 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11799 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11800 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 11801 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 11802 then
	sram_write <= x"005A0000";
end if;
if first_state_sram_input_id = 11803 then
	sram_write <= x"03BA0008";
end if;
if first_state_sram_input_id = 11804 then
	sram_write <= x"C4240004";
end if;
if first_state_sram_input_id = 11805 then
	sram_write <= x"C03C0024";
end if;
if first_state_sram_input_id = 11806 then
	sram_write <= x"C4240000";
end if;
if first_state_sram_input_id = 11807 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 11808 then
	sram_write <= x"C05C0020";
end if;
if first_state_sram_input_id = 11809 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 11810 then
	sram_write <= x"C09C0008";
end if;
if first_state_sram_input_id = 11811 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 11812 then
	sram_write <= x"06240001";
end if;
if first_state_sram_input_id = 11813 then
	sram_write <= x"8620B91C";
end if;
if first_state_sram_input_id = 11814 then
	sram_write <= x"02400003";
end if;
if first_state_sram_input_id = 11815 then
	sram_write <= x"C83C0000";
end if;
if first_state_sram_input_id = 11816 then
	sram_write <= x"C43C0028";
end if;
if first_state_sram_input_id = 11817 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11818 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 11819 then
	sram_write <= x"03DC0034";
end if;
if first_state_sram_input_id = 11820 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11821 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11822 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 11823 then
	sram_write <= x"07DC0034";
end if;
if first_state_sram_input_id = 11824 then
	sram_write <= x"00420000";
end if;
if first_state_sram_input_id = 11825 then
	sram_write <= x"C03C0010";
end if;
if first_state_sram_input_id = 11826 then
	sram_write <= x"C0220000";
end if;
if first_state_sram_input_id = 11827 then
	sram_write <= x"C45C002C";
end if;
if first_state_sram_input_id = 11828 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11829 then
	sram_write <= x"03DC0038";
end if;
if first_state_sram_input_id = 11830 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11831 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11832 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 11833 then
	sram_write <= x"07DC0038";
end if;
if first_state_sram_input_id = 11834 then
	sram_write <= x"005A0000";
end if;
if first_state_sram_input_id = 11835 then
	sram_write <= x"03BA0008";
end if;
if first_state_sram_input_id = 11836 then
	sram_write <= x"C4240004";
end if;
if first_state_sram_input_id = 11837 then
	sram_write <= x"C03C002C";
end if;
if first_state_sram_input_id = 11838 then
	sram_write <= x"C4240000";
end if;
if first_state_sram_input_id = 11839 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 11840 then
	sram_write <= x"C05C0028";
end if;
if first_state_sram_input_id = 11841 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 11842 then
	sram_write <= x"C09C0008";
end if;
if first_state_sram_input_id = 11843 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 11844 then
	sram_write <= x"06440001";
end if;
if first_state_sram_input_id = 11845 then
	sram_write <= x"00280000";
end if;
if first_state_sram_input_id = 11846 then
	sram_write <= x"8200B6FC";
end if;
if first_state_sram_input_id = 11847 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 11848 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 11849 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 11850 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 11851 then
	sram_write <= x"8620BD0C";
end if;
if first_state_sram_input_id = 11852 then
	sram_write <= x"02400354";
end if;
if first_state_sram_input_id = 11853 then
	sram_write <= x"02600078";
end if;
if first_state_sram_input_id = 11854 then
	sram_write <= x"02800003";
end if;
if first_state_sram_input_id = 11855 then
	sram_write <= x"40200000";
end if;
if first_state_sram_input_id = 11856 then
	sram_write <= x"CC3C0000";
end if;
if first_state_sram_input_id = 11857 then
	sram_write <= x"C45C0008";
end if;
if first_state_sram_input_id = 11858 then
	sram_write <= x"C43C000C";
end if;
if first_state_sram_input_id = 11859 then
	sram_write <= x"C47C0010";
end if;
if first_state_sram_input_id = 11860 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11861 then
	sram_write <= x"00280000";
end if;
if first_state_sram_input_id = 11862 then
	sram_write <= x"03DC001C";
end if;
if first_state_sram_input_id = 11863 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11864 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11865 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 11866 then
	sram_write <= x"07DC001C";
end if;
if first_state_sram_input_id = 11867 then
	sram_write <= x"00420000";
end if;
if first_state_sram_input_id = 11868 then
	sram_write <= x"022000C4";
end if;
if first_state_sram_input_id = 11869 then
	sram_write <= x"C0620000";
end if;
if first_state_sram_input_id = 11870 then
	sram_write <= x"C43C0014";
end if;
if first_state_sram_input_id = 11871 then
	sram_write <= x"C45C0018";
end if;
if first_state_sram_input_id = 11872 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11873 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 11874 then
	sram_write <= x"03DC0024";
end if;
if first_state_sram_input_id = 11875 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11876 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11877 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 11878 then
	sram_write <= x"07DC0024";
end if;
if first_state_sram_input_id = 11879 then
	sram_write <= x"005A0000";
end if;
if first_state_sram_input_id = 11880 then
	sram_write <= x"03BA0008";
end if;
if first_state_sram_input_id = 11881 then
	sram_write <= x"C4240004";
end if;
if first_state_sram_input_id = 11882 then
	sram_write <= x"C03C0018";
end if;
if first_state_sram_input_id = 11883 then
	sram_write <= x"C4240000";
end if;
if first_state_sram_input_id = 11884 then
	sram_write <= x"C03C0010";
end if;
if first_state_sram_input_id = 11885 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11886 then
	sram_write <= x"03DC0024";
end if;
if first_state_sram_input_id = 11887 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11888 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11889 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 11890 then
	sram_write <= x"07DC0024";
end if;
if first_state_sram_input_id = 11891 then
	sram_write <= x"C05C000C";
end if;
if first_state_sram_input_id = 11892 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 11893 then
	sram_write <= x"C09C0008";
end if;
if first_state_sram_input_id = 11894 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 11895 then
	sram_write <= x"02600003";
end if;
if first_state_sram_input_id = 11896 then
	sram_write <= x"C83C0000";
end if;
if first_state_sram_input_id = 11897 then
	sram_write <= x"C43C001C";
end if;
if first_state_sram_input_id = 11898 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11899 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 11900 then
	sram_write <= x"03DC0028";
end if;
if first_state_sram_input_id = 11901 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11902 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11903 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 11904 then
	sram_write <= x"07DC0028";
end if;
if first_state_sram_input_id = 11905 then
	sram_write <= x"00420000";
end if;
if first_state_sram_input_id = 11906 then
	sram_write <= x"C03C0014";
end if;
if first_state_sram_input_id = 11907 then
	sram_write <= x"C0620000";
end if;
if first_state_sram_input_id = 11908 then
	sram_write <= x"C45C0020";
end if;
if first_state_sram_input_id = 11909 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11910 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 11911 then
	sram_write <= x"03DC002C";
end if;
if first_state_sram_input_id = 11912 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11913 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11914 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 11915 then
	sram_write <= x"07DC002C";
end if;
if first_state_sram_input_id = 11916 then
	sram_write <= x"005A0000";
end if;
if first_state_sram_input_id = 11917 then
	sram_write <= x"03BA0008";
end if;
if first_state_sram_input_id = 11918 then
	sram_write <= x"C4240004";
end if;
if first_state_sram_input_id = 11919 then
	sram_write <= x"C03C0020";
end if;
if first_state_sram_input_id = 11920 then
	sram_write <= x"C4240000";
end if;
if first_state_sram_input_id = 11921 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 11922 then
	sram_write <= x"C05C001C";
end if;
if first_state_sram_input_id = 11923 then
	sram_write <= x"C42401D8";
end if;
if first_state_sram_input_id = 11924 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 11925 then
	sram_write <= x"C83C0000";
end if;
if first_state_sram_input_id = 11926 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11927 then
	sram_write <= x"03DC002C";
end if;
if first_state_sram_input_id = 11928 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11929 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11930 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 11931 then
	sram_write <= x"07DC002C";
end if;
if first_state_sram_input_id = 11932 then
	sram_write <= x"00420000";
end if;
if first_state_sram_input_id = 11933 then
	sram_write <= x"C03C0014";
end if;
if first_state_sram_input_id = 11934 then
	sram_write <= x"C0620000";
end if;
if first_state_sram_input_id = 11935 then
	sram_write <= x"C45C0024";
end if;
if first_state_sram_input_id = 11936 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11937 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 11938 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 11939 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11940 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11941 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 11942 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 11943 then
	sram_write <= x"005A0000";
end if;
if first_state_sram_input_id = 11944 then
	sram_write <= x"03BA0008";
end if;
if first_state_sram_input_id = 11945 then
	sram_write <= x"C4240004";
end if;
if first_state_sram_input_id = 11946 then
	sram_write <= x"C03C0024";
end if;
if first_state_sram_input_id = 11947 then
	sram_write <= x"C4240000";
end if;
if first_state_sram_input_id = 11948 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 11949 then
	sram_write <= x"C05C001C";
end if;
if first_state_sram_input_id = 11950 then
	sram_write <= x"C42401D4";
end if;
if first_state_sram_input_id = 11951 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 11952 then
	sram_write <= x"C83C0000";
end if;
if first_state_sram_input_id = 11953 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11954 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 11955 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11956 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11957 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 11958 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 11959 then
	sram_write <= x"00420000";
end if;
if first_state_sram_input_id = 11960 then
	sram_write <= x"C03C0014";
end if;
if first_state_sram_input_id = 11961 then
	sram_write <= x"C0620000";
end if;
if first_state_sram_input_id = 11962 then
	sram_write <= x"C45C0028";
end if;
if first_state_sram_input_id = 11963 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11964 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 11965 then
	sram_write <= x"03DC0034";
end if;
if first_state_sram_input_id = 11966 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11967 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11968 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 11969 then
	sram_write <= x"07DC0034";
end if;
if first_state_sram_input_id = 11970 then
	sram_write <= x"005A0000";
end if;
if first_state_sram_input_id = 11971 then
	sram_write <= x"03BA0008";
end if;
if first_state_sram_input_id = 11972 then
	sram_write <= x"C4240004";
end if;
if first_state_sram_input_id = 11973 then
	sram_write <= x"C03C0028";
end if;
if first_state_sram_input_id = 11974 then
	sram_write <= x"C4240000";
end if;
if first_state_sram_input_id = 11975 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 11976 then
	sram_write <= x"C05C001C";
end if;
if first_state_sram_input_id = 11977 then
	sram_write <= x"C42401D0";
end if;
if first_state_sram_input_id = 11978 then
	sram_write <= x"02200073";
end if;
if first_state_sram_input_id = 11979 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11980 then
	sram_write <= x"01240000";
end if;
if first_state_sram_input_id = 11981 then
	sram_write <= x"00420000";
end if;
if first_state_sram_input_id = 11982 then
	sram_write <= x"00320000";
end if;
if first_state_sram_input_id = 11983 then
	sram_write <= x"03DC0034";
end if;
if first_state_sram_input_id = 11984 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 11985 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 11986 then
	sram_write <= x"8200B6FC";
end if;
if first_state_sram_input_id = 11987 then
	sram_write <= x"07DC0034";
end if;
if first_state_sram_input_id = 11988 then
	sram_write <= x"C03C000C";
end if;
if first_state_sram_input_id = 11989 then
	sram_write <= x"06220001";
end if;
if first_state_sram_input_id = 11990 then
	sram_write <= x"8620BD08";
end if;
if first_state_sram_input_id = 11991 then
	sram_write <= x"02400078";
end if;
if first_state_sram_input_id = 11992 then
	sram_write <= x"02600003";
end if;
if first_state_sram_input_id = 11993 then
	sram_write <= x"C83C0000";
end if;
if first_state_sram_input_id = 11994 then
	sram_write <= x"C43C002C";
end if;
if first_state_sram_input_id = 11995 then
	sram_write <= x"C45C0030";
end if;
if first_state_sram_input_id = 11996 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 11997 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 11998 then
	sram_write <= x"03DC003C";
end if;
if first_state_sram_input_id = 11999 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12000 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12001 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 12002 then
	sram_write <= x"07DC003C";
end if;
if first_state_sram_input_id = 12003 then
	sram_write <= x"00420000";
end if;
if first_state_sram_input_id = 12004 then
	sram_write <= x"C03C0014";
end if;
if first_state_sram_input_id = 12005 then
	sram_write <= x"C0620000";
end if;
if first_state_sram_input_id = 12006 then
	sram_write <= x"C45C0034";
end if;
if first_state_sram_input_id = 12007 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12008 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 12009 then
	sram_write <= x"03DC0040";
end if;
if first_state_sram_input_id = 12010 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12011 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12012 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 12013 then
	sram_write <= x"07DC0040";
end if;
if first_state_sram_input_id = 12014 then
	sram_write <= x"005A0000";
end if;
if first_state_sram_input_id = 12015 then
	sram_write <= x"03BA0008";
end if;
if first_state_sram_input_id = 12016 then
	sram_write <= x"C4240004";
end if;
if first_state_sram_input_id = 12017 then
	sram_write <= x"C03C0034";
end if;
if first_state_sram_input_id = 12018 then
	sram_write <= x"C4240000";
end if;
if first_state_sram_input_id = 12019 then
	sram_write <= x"C03C0030";
end if;
if first_state_sram_input_id = 12020 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12021 then
	sram_write <= x"03DC0040";
end if;
if first_state_sram_input_id = 12022 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12023 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12024 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 12025 then
	sram_write <= x"07DC0040";
end if;
if first_state_sram_input_id = 12026 then
	sram_write <= x"C05C002C";
end if;
if first_state_sram_input_id = 12027 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 12028 then
	sram_write <= x"C09C0008";
end if;
if first_state_sram_input_id = 12029 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 12030 then
	sram_write <= x"02600003";
end if;
if first_state_sram_input_id = 12031 then
	sram_write <= x"C83C0000";
end if;
if first_state_sram_input_id = 12032 then
	sram_write <= x"C43C0038";
end if;
if first_state_sram_input_id = 12033 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12034 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 12035 then
	sram_write <= x"03DC0044";
end if;
if first_state_sram_input_id = 12036 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12037 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12038 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 12039 then
	sram_write <= x"07DC0044";
end if;
if first_state_sram_input_id = 12040 then
	sram_write <= x"00420000";
end if;
if first_state_sram_input_id = 12041 then
	sram_write <= x"C03C0014";
end if;
if first_state_sram_input_id = 12042 then
	sram_write <= x"C0620000";
end if;
if first_state_sram_input_id = 12043 then
	sram_write <= x"C45C003C";
end if;
if first_state_sram_input_id = 12044 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12045 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 12046 then
	sram_write <= x"03DC0048";
end if;
if first_state_sram_input_id = 12047 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12048 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12049 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 12050 then
	sram_write <= x"07DC0048";
end if;
if first_state_sram_input_id = 12051 then
	sram_write <= x"005A0000";
end if;
if first_state_sram_input_id = 12052 then
	sram_write <= x"03BA0008";
end if;
if first_state_sram_input_id = 12053 then
	sram_write <= x"C4240004";
end if;
if first_state_sram_input_id = 12054 then
	sram_write <= x"C03C003C";
end if;
if first_state_sram_input_id = 12055 then
	sram_write <= x"C4240000";
end if;
if first_state_sram_input_id = 12056 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 12057 then
	sram_write <= x"C05C0038";
end if;
if first_state_sram_input_id = 12058 then
	sram_write <= x"C42401D8";
end if;
if first_state_sram_input_id = 12059 then
	sram_write <= x"02200003";
end if;
if first_state_sram_input_id = 12060 then
	sram_write <= x"C83C0000";
end if;
if first_state_sram_input_id = 12061 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12062 then
	sram_write <= x"03DC0048";
end if;
if first_state_sram_input_id = 12063 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12064 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12065 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 12066 then
	sram_write <= x"07DC0048";
end if;
if first_state_sram_input_id = 12067 then
	sram_write <= x"00420000";
end if;
if first_state_sram_input_id = 12068 then
	sram_write <= x"C03C0014";
end if;
if first_state_sram_input_id = 12069 then
	sram_write <= x"C0220000";
end if;
if first_state_sram_input_id = 12070 then
	sram_write <= x"C45C0040";
end if;
if first_state_sram_input_id = 12071 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12072 then
	sram_write <= x"03DC004C";
end if;
if first_state_sram_input_id = 12073 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12074 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12075 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 12076 then
	sram_write <= x"07DC004C";
end if;
if first_state_sram_input_id = 12077 then
	sram_write <= x"005A0000";
end if;
if first_state_sram_input_id = 12078 then
	sram_write <= x"03BA0008";
end if;
if first_state_sram_input_id = 12079 then
	sram_write <= x"C4240004";
end if;
if first_state_sram_input_id = 12080 then
	sram_write <= x"C03C0040";
end if;
if first_state_sram_input_id = 12081 then
	sram_write <= x"C4240000";
end if;
if first_state_sram_input_id = 12082 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 12083 then
	sram_write <= x"C05C0038";
end if;
if first_state_sram_input_id = 12084 then
	sram_write <= x"C42401D4";
end if;
if first_state_sram_input_id = 12085 then
	sram_write <= x"02200074";
end if;
if first_state_sram_input_id = 12086 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12087 then
	sram_write <= x"01240000";
end if;
if first_state_sram_input_id = 12088 then
	sram_write <= x"00420000";
end if;
if first_state_sram_input_id = 12089 then
	sram_write <= x"00320000";
end if;
if first_state_sram_input_id = 12090 then
	sram_write <= x"03DC004C";
end if;
if first_state_sram_input_id = 12091 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12092 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12093 then
	sram_write <= x"8200B6FC";
end if;
if first_state_sram_input_id = 12094 then
	sram_write <= x"07DC004C";
end if;
if first_state_sram_input_id = 12095 then
	sram_write <= x"C03C002C";
end if;
if first_state_sram_input_id = 12096 then
	sram_write <= x"06220001";
end if;
if first_state_sram_input_id = 12097 then
	sram_write <= x"8200B92C";
end if;
if first_state_sram_input_id = 12098 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 12099 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 12100 then
	sram_write <= x"8640C710";
end if;
if first_state_sram_input_id = 12101 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 12102 then
	sram_write <= x"D0626000";
end if;
if first_state_sram_input_id = 12103 then
	sram_write <= x"028000C4";
end if;
if first_state_sram_input_id = 12104 then
	sram_write <= x"C0A80000";
end if;
if first_state_sram_input_id = 12105 then
	sram_write <= x"06AA0001";
end if;
if first_state_sram_input_id = 12106 then
	sram_write <= x"C49C0000";
end if;
if first_state_sram_input_id = 12107 then
	sram_write <= x"C43C0004";
end if;
if first_state_sram_input_id = 12108 then
	sram_write <= x"C45C0008";
end if;
if first_state_sram_input_id = 12109 then
	sram_write <= x"86A0BF18";
end if;
if first_state_sram_input_id = 12110 then
	sram_write <= x"02C000C8";
end if;
if first_state_sram_input_id = 12111 then
	sram_write <= x"22EA0220";
end if;
if first_state_sram_input_id = 12112 then
	sram_write <= x"D0ECE000";
end if;
if first_state_sram_input_id = 12113 then
	sram_write <= x"C1060004";
end if;
if first_state_sram_input_id = 12114 then
	sram_write <= x"C1260000";
end if;
if first_state_sram_input_id = 12115 then
	sram_write <= x"C14E0004";
end if;
if first_state_sram_input_id = 12116 then
	sram_write <= x"02800001";
end if;
if first_state_sram_input_id = 12117 then
	sram_write <= x"C47C000C";
end if;
if first_state_sram_input_id = 12118 then
	sram_write <= x"C4DC0010";
end if;
if first_state_sram_input_id = 12119 then
	sram_write <= x"8348BDE0";
end if;
if first_state_sram_input_id = 12120 then
	sram_write <= x"02800002";
end if;
if first_state_sram_input_id = 12121 then
	sram_write <= x"8348BDA4";
end if;
if first_state_sram_input_id = 12122 then
	sram_write <= x"C51C0014";
end if;
if first_state_sram_input_id = 12123 then
	sram_write <= x"C4BC0018";
end if;
if first_state_sram_input_id = 12124 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12125 then
	sram_write <= x"004E0000";
end if;
if first_state_sram_input_id = 12126 then
	sram_write <= x"00320000";
end if;
if first_state_sram_input_id = 12127 then
	sram_write <= x"03DC0024";
end if;
if first_state_sram_input_id = 12128 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12129 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12130 then
	sram_write <= x"8200400C";
end if;
if first_state_sram_input_id = 12131 then
	sram_write <= x"07DC0024";
end if;
if first_state_sram_input_id = 12132 then
	sram_write <= x"C05C0018";
end if;
if first_state_sram_input_id = 12133 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 12134 then
	sram_write <= x"C09C0014";
end if;
if first_state_sram_input_id = 12135 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 12136 then
	sram_write <= x"8200BDDC";
end if;
if first_state_sram_input_id = 12137 then
	sram_write <= x"C51C0014";
end if;
if first_state_sram_input_id = 12138 then
	sram_write <= x"C4BC0018";
end if;
if first_state_sram_input_id = 12139 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12140 then
	sram_write <= x"004E0000";
end if;
if first_state_sram_input_id = 12141 then
	sram_write <= x"00320000";
end if;
if first_state_sram_input_id = 12142 then
	sram_write <= x"03DC0024";
end if;
if first_state_sram_input_id = 12143 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12144 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12145 then
	sram_write <= x"82003E98";
end if;
if first_state_sram_input_id = 12146 then
	sram_write <= x"07DC0024";
end if;
if first_state_sram_input_id = 12147 then
	sram_write <= x"C05C0018";
end if;
if first_state_sram_input_id = 12148 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 12149 then
	sram_write <= x"C09C0014";
end if;
if first_state_sram_input_id = 12150 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 12151 then
	sram_write <= x"8200BE18";
end if;
if first_state_sram_input_id = 12152 then
	sram_write <= x"C51C0014";
end if;
if first_state_sram_input_id = 12153 then
	sram_write <= x"C4BC0018";
end if;
if first_state_sram_input_id = 12154 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12155 then
	sram_write <= x"004E0000";
end if;
if first_state_sram_input_id = 12156 then
	sram_write <= x"00320000";
end if;
if first_state_sram_input_id = 12157 then
	sram_write <= x"03DC0024";
end if;
if first_state_sram_input_id = 12158 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12159 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12160 then
	sram_write <= x"82003CC4";
end if;
if first_state_sram_input_id = 12161 then
	sram_write <= x"07DC0024";
end if;
if first_state_sram_input_id = 12162 then
	sram_write <= x"C05C0018";
end if;
if first_state_sram_input_id = 12163 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 12164 then
	sram_write <= x"C09C0014";
end if;
if first_state_sram_input_id = 12165 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 12166 then
	sram_write <= x"06240001";
end if;
if first_state_sram_input_id = 12167 then
	sram_write <= x"8620BF14";
end if;
if first_state_sram_input_id = 12168 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 12169 then
	sram_write <= x"C07C0010";
end if;
if first_state_sram_input_id = 12170 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 12171 then
	sram_write <= x"C07C000C";
end if;
if first_state_sram_input_id = 12172 then
	sram_write <= x"C0860004";
end if;
if first_state_sram_input_id = 12173 then
	sram_write <= x"C0A60000";
end if;
if first_state_sram_input_id = 12174 then
	sram_write <= x"C0C40004";
end if;
if first_state_sram_input_id = 12175 then
	sram_write <= x"02E00001";
end if;
if first_state_sram_input_id = 12176 then
	sram_write <= x"82CEBEBC";
end if;
if first_state_sram_input_id = 12177 then
	sram_write <= x"02E00002";
end if;
if first_state_sram_input_id = 12178 then
	sram_write <= x"82CEBE84";
end if;
if first_state_sram_input_id = 12179 then
	sram_write <= x"C49C001C";
end if;
if first_state_sram_input_id = 12180 then
	sram_write <= x"C43C0020";
end if;
if first_state_sram_input_id = 12181 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12182 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 12183 then
	sram_write <= x"03DC002C";
end if;
if first_state_sram_input_id = 12184 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12185 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12186 then
	sram_write <= x"8200400C";
end if;
if first_state_sram_input_id = 12187 then
	sram_write <= x"07DC002C";
end if;
if first_state_sram_input_id = 12188 then
	sram_write <= x"C05C0020";
end if;
if first_state_sram_input_id = 12189 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 12190 then
	sram_write <= x"C09C001C";
end if;
if first_state_sram_input_id = 12191 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 12192 then
	sram_write <= x"8200BEB8";
end if;
if first_state_sram_input_id = 12193 then
	sram_write <= x"C49C001C";
end if;
if first_state_sram_input_id = 12194 then
	sram_write <= x"C43C0020";
end if;
if first_state_sram_input_id = 12195 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12196 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 12197 then
	sram_write <= x"03DC002C";
end if;
if first_state_sram_input_id = 12198 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12199 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12200 then
	sram_write <= x"82003E98";
end if;
if first_state_sram_input_id = 12201 then
	sram_write <= x"07DC002C";
end if;
if first_state_sram_input_id = 12202 then
	sram_write <= x"C05C0020";
end if;
if first_state_sram_input_id = 12203 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 12204 then
	sram_write <= x"C09C001C";
end if;
if first_state_sram_input_id = 12205 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 12206 then
	sram_write <= x"8200BEF0";
end if;
if first_state_sram_input_id = 12207 then
	sram_write <= x"C49C001C";
end if;
if first_state_sram_input_id = 12208 then
	sram_write <= x"C43C0020";
end if;
if first_state_sram_input_id = 12209 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12210 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 12211 then
	sram_write <= x"03DC002C";
end if;
if first_state_sram_input_id = 12212 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12213 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12214 then
	sram_write <= x"82003CC4";
end if;
if first_state_sram_input_id = 12215 then
	sram_write <= x"07DC002C";
end if;
if first_state_sram_input_id = 12216 then
	sram_write <= x"C05C0020";
end if;
if first_state_sram_input_id = 12217 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 12218 then
	sram_write <= x"C09C001C";
end if;
if first_state_sram_input_id = 12219 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 12220 then
	sram_write <= x"06440001";
end if;
if first_state_sram_input_id = 12221 then
	sram_write <= x"C03C000C";
end if;
if first_state_sram_input_id = 12222 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12223 then
	sram_write <= x"03DC002C";
end if;
if first_state_sram_input_id = 12224 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12225 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12226 then
	sram_write <= x"820042A4";
end if;
if first_state_sram_input_id = 12227 then
	sram_write <= x"07DC002C";
end if;
if first_state_sram_input_id = 12228 then
	sram_write <= x"8200BF14";
end if;
if first_state_sram_input_id = 12229 then
	sram_write <= x"8200BF18";
end if;
if first_state_sram_input_id = 12230 then
	sram_write <= x"C03C0008";
end if;
if first_state_sram_input_id = 12231 then
	sram_write <= x"06220001";
end if;
if first_state_sram_input_id = 12232 then
	sram_write <= x"8620C70C";
end if;
if first_state_sram_input_id = 12233 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 12234 then
	sram_write <= x"C07C0004";
end if;
if first_state_sram_input_id = 12235 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 12236 then
	sram_write <= x"C09C0000";
end if;
if first_state_sram_input_id = 12237 then
	sram_write <= x"C0A80000";
end if;
if first_state_sram_input_id = 12238 then
	sram_write <= x"06AA0001";
end if;
if first_state_sram_input_id = 12239 then
	sram_write <= x"C43C0024";
end if;
if first_state_sram_input_id = 12240 then
	sram_write <= x"86A0C200";
end if;
if first_state_sram_input_id = 12241 then
	sram_write <= x"02C000C8";
end if;
if first_state_sram_input_id = 12242 then
	sram_write <= x"22EA0220";
end if;
if first_state_sram_input_id = 12243 then
	sram_write <= x"D0ECE000";
end if;
if first_state_sram_input_id = 12244 then
	sram_write <= x"C1040004";
end if;
if first_state_sram_input_id = 12245 then
	sram_write <= x"C1240000";
end if;
if first_state_sram_input_id = 12246 then
	sram_write <= x"C14E0004";
end if;
if first_state_sram_input_id = 12247 then
	sram_write <= x"02800001";
end if;
if first_state_sram_input_id = 12248 then
	sram_write <= x"C45C0028";
end if;
if first_state_sram_input_id = 12249 then
	sram_write <= x"C4DC002C";
end if;
if first_state_sram_input_id = 12250 then
	sram_write <= x"8348BFEC";
end if;
if first_state_sram_input_id = 12251 then
	sram_write <= x"02800002";
end if;
if first_state_sram_input_id = 12252 then
	sram_write <= x"8348BFB0";
end if;
if first_state_sram_input_id = 12253 then
	sram_write <= x"C51C0030";
end if;
if first_state_sram_input_id = 12254 then
	sram_write <= x"C4BC0034";
end if;
if first_state_sram_input_id = 12255 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12256 then
	sram_write <= x"004E0000";
end if;
if first_state_sram_input_id = 12257 then
	sram_write <= x"00320000";
end if;
if first_state_sram_input_id = 12258 then
	sram_write <= x"03DC0040";
end if;
if first_state_sram_input_id = 12259 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12260 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12261 then
	sram_write <= x"8200400C";
end if;
if first_state_sram_input_id = 12262 then
	sram_write <= x"07DC0040";
end if;
if first_state_sram_input_id = 12263 then
	sram_write <= x"C05C0034";
end if;
if first_state_sram_input_id = 12264 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 12265 then
	sram_write <= x"C09C0030";
end if;
if first_state_sram_input_id = 12266 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 12267 then
	sram_write <= x"8200BFE8";
end if;
if first_state_sram_input_id = 12268 then
	sram_write <= x"C51C0030";
end if;
if first_state_sram_input_id = 12269 then
	sram_write <= x"C4BC0034";
end if;
if first_state_sram_input_id = 12270 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12271 then
	sram_write <= x"004E0000";
end if;
if first_state_sram_input_id = 12272 then
	sram_write <= x"00320000";
end if;
if first_state_sram_input_id = 12273 then
	sram_write <= x"03DC0040";
end if;
if first_state_sram_input_id = 12274 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12275 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12276 then
	sram_write <= x"82003E98";
end if;
if first_state_sram_input_id = 12277 then
	sram_write <= x"07DC0040";
end if;
if first_state_sram_input_id = 12278 then
	sram_write <= x"C05C0034";
end if;
if first_state_sram_input_id = 12279 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 12280 then
	sram_write <= x"C09C0030";
end if;
if first_state_sram_input_id = 12281 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 12282 then
	sram_write <= x"8200C024";
end if;
if first_state_sram_input_id = 12283 then
	sram_write <= x"C51C0030";
end if;
if first_state_sram_input_id = 12284 then
	sram_write <= x"C4BC0034";
end if;
if first_state_sram_input_id = 12285 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12286 then
	sram_write <= x"004E0000";
end if;
if first_state_sram_input_id = 12287 then
	sram_write <= x"00320000";
end if;
if first_state_sram_input_id = 12288 then
	sram_write <= x"03DC0040";
end if;
if first_state_sram_input_id = 12289 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12290 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12291 then
	sram_write <= x"82003CC4";
end if;
if first_state_sram_input_id = 12292 then
	sram_write <= x"07DC0040";
end if;
if first_state_sram_input_id = 12293 then
	sram_write <= x"C05C0034";
end if;
if first_state_sram_input_id = 12294 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 12295 then
	sram_write <= x"C09C0030";
end if;
if first_state_sram_input_id = 12296 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 12297 then
	sram_write <= x"06240001";
end if;
if first_state_sram_input_id = 12298 then
	sram_write <= x"8620C1FC";
end if;
if first_state_sram_input_id = 12299 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 12300 then
	sram_write <= x"C07C002C";
end if;
if first_state_sram_input_id = 12301 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 12302 then
	sram_write <= x"C09C0028";
end if;
if first_state_sram_input_id = 12303 then
	sram_write <= x"C0A80004";
end if;
if first_state_sram_input_id = 12304 then
	sram_write <= x"C0C80000";
end if;
if first_state_sram_input_id = 12305 then
	sram_write <= x"C0E40004";
end if;
if first_state_sram_input_id = 12306 then
	sram_write <= x"03000001";
end if;
if first_state_sram_input_id = 12307 then
	sram_write <= x"82F0C0C8";
end if;
if first_state_sram_input_id = 12308 then
	sram_write <= x"03000002";
end if;
if first_state_sram_input_id = 12309 then
	sram_write <= x"82F0C090";
end if;
if first_state_sram_input_id = 12310 then
	sram_write <= x"C4BC0038";
end if;
if first_state_sram_input_id = 12311 then
	sram_write <= x"C43C003C";
end if;
if first_state_sram_input_id = 12312 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12313 then
	sram_write <= x"002C0000";
end if;
if first_state_sram_input_id = 12314 then
	sram_write <= x"03DC0048";
end if;
if first_state_sram_input_id = 12315 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12316 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12317 then
	sram_write <= x"8200400C";
end if;
if first_state_sram_input_id = 12318 then
	sram_write <= x"07DC0048";
end if;
if first_state_sram_input_id = 12319 then
	sram_write <= x"C05C003C";
end if;
if first_state_sram_input_id = 12320 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 12321 then
	sram_write <= x"C09C0038";
end if;
if first_state_sram_input_id = 12322 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 12323 then
	sram_write <= x"8200C0C4";
end if;
if first_state_sram_input_id = 12324 then
	sram_write <= x"C4BC0038";
end if;
if first_state_sram_input_id = 12325 then
	sram_write <= x"C43C003C";
end if;
if first_state_sram_input_id = 12326 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12327 then
	sram_write <= x"002C0000";
end if;
if first_state_sram_input_id = 12328 then
	sram_write <= x"03DC0048";
end if;
if first_state_sram_input_id = 12329 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12330 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12331 then
	sram_write <= x"82003E98";
end if;
if first_state_sram_input_id = 12332 then
	sram_write <= x"07DC0048";
end if;
if first_state_sram_input_id = 12333 then
	sram_write <= x"C05C003C";
end if;
if first_state_sram_input_id = 12334 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 12335 then
	sram_write <= x"C09C0038";
end if;
if first_state_sram_input_id = 12336 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 12337 then
	sram_write <= x"8200C0FC";
end if;
if first_state_sram_input_id = 12338 then
	sram_write <= x"C4BC0038";
end if;
if first_state_sram_input_id = 12339 then
	sram_write <= x"C43C003C";
end if;
if first_state_sram_input_id = 12340 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12341 then
	sram_write <= x"002C0000";
end if;
if first_state_sram_input_id = 12342 then
	sram_write <= x"03DC0048";
end if;
if first_state_sram_input_id = 12343 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12344 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12345 then
	sram_write <= x"82003CC4";
end if;
if first_state_sram_input_id = 12346 then
	sram_write <= x"07DC0048";
end if;
if first_state_sram_input_id = 12347 then
	sram_write <= x"C05C003C";
end if;
if first_state_sram_input_id = 12348 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 12349 then
	sram_write <= x"C09C0038";
end if;
if first_state_sram_input_id = 12350 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 12351 then
	sram_write <= x"06240001";
end if;
if first_state_sram_input_id = 12352 then
	sram_write <= x"8620C1F8";
end if;
if first_state_sram_input_id = 12353 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 12354 then
	sram_write <= x"C07C002C";
end if;
if first_state_sram_input_id = 12355 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 12356 then
	sram_write <= x"C07C0028";
end if;
if first_state_sram_input_id = 12357 then
	sram_write <= x"C0860004";
end if;
if first_state_sram_input_id = 12358 then
	sram_write <= x"C0A60000";
end if;
if first_state_sram_input_id = 12359 then
	sram_write <= x"C0C40004";
end if;
if first_state_sram_input_id = 12360 then
	sram_write <= x"02E00001";
end if;
if first_state_sram_input_id = 12361 then
	sram_write <= x"82CEC1A0";
end if;
if first_state_sram_input_id = 12362 then
	sram_write <= x"02E00002";
end if;
if first_state_sram_input_id = 12363 then
	sram_write <= x"82CEC168";
end if;
if first_state_sram_input_id = 12364 then
	sram_write <= x"C49C0040";
end if;
if first_state_sram_input_id = 12365 then
	sram_write <= x"C43C0044";
end if;
if first_state_sram_input_id = 12366 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12367 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 12368 then
	sram_write <= x"03DC0050";
end if;
if first_state_sram_input_id = 12369 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12370 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12371 then
	sram_write <= x"8200400C";
end if;
if first_state_sram_input_id = 12372 then
	sram_write <= x"07DC0050";
end if;
if first_state_sram_input_id = 12373 then
	sram_write <= x"C05C0044";
end if;
if first_state_sram_input_id = 12374 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 12375 then
	sram_write <= x"C09C0040";
end if;
if first_state_sram_input_id = 12376 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 12377 then
	sram_write <= x"8200C19C";
end if;
if first_state_sram_input_id = 12378 then
	sram_write <= x"C49C0040";
end if;
if first_state_sram_input_id = 12379 then
	sram_write <= x"C43C0044";
end if;
if first_state_sram_input_id = 12380 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12381 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 12382 then
	sram_write <= x"03DC0050";
end if;
if first_state_sram_input_id = 12383 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12384 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12385 then
	sram_write <= x"82003E98";
end if;
if first_state_sram_input_id = 12386 then
	sram_write <= x"07DC0050";
end if;
if first_state_sram_input_id = 12387 then
	sram_write <= x"C05C0044";
end if;
if first_state_sram_input_id = 12388 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 12389 then
	sram_write <= x"C09C0040";
end if;
if first_state_sram_input_id = 12390 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 12391 then
	sram_write <= x"8200C1D4";
end if;
if first_state_sram_input_id = 12392 then
	sram_write <= x"C49C0040";
end if;
if first_state_sram_input_id = 12393 then
	sram_write <= x"C43C0044";
end if;
if first_state_sram_input_id = 12394 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12395 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 12396 then
	sram_write <= x"03DC0050";
end if;
if first_state_sram_input_id = 12397 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12398 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12399 then
	sram_write <= x"82003CC4";
end if;
if first_state_sram_input_id = 12400 then
	sram_write <= x"07DC0050";
end if;
if first_state_sram_input_id = 12401 then
	sram_write <= x"C05C0044";
end if;
if first_state_sram_input_id = 12402 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 12403 then
	sram_write <= x"C09C0040";
end if;
if first_state_sram_input_id = 12404 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 12405 then
	sram_write <= x"06440001";
end if;
if first_state_sram_input_id = 12406 then
	sram_write <= x"C03C0028";
end if;
if first_state_sram_input_id = 12407 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12408 then
	sram_write <= x"03DC0050";
end if;
if first_state_sram_input_id = 12409 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12410 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12411 then
	sram_write <= x"820042A4";
end if;
if first_state_sram_input_id = 12412 then
	sram_write <= x"07DC0050";
end if;
if first_state_sram_input_id = 12413 then
	sram_write <= x"8200C1F8";
end if;
if first_state_sram_input_id = 12414 then
	sram_write <= x"8200C1FC";
end if;
if first_state_sram_input_id = 12415 then
	sram_write <= x"8200C200";
end if;
if first_state_sram_input_id = 12416 then
	sram_write <= x"C03C0024";
end if;
if first_state_sram_input_id = 12417 then
	sram_write <= x"06220001";
end if;
if first_state_sram_input_id = 12418 then
	sram_write <= x"8620C708";
end if;
if first_state_sram_input_id = 12419 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 12420 then
	sram_write <= x"C07C0004";
end if;
if first_state_sram_input_id = 12421 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 12422 then
	sram_write <= x"C09C0000";
end if;
if first_state_sram_input_id = 12423 then
	sram_write <= x"C0A80000";
end if;
if first_state_sram_input_id = 12424 then
	sram_write <= x"06AA0001";
end if;
if first_state_sram_input_id = 12425 then
	sram_write <= x"C43C0048";
end if;
if first_state_sram_input_id = 12426 then
	sram_write <= x"86A0C40C";
end if;
if first_state_sram_input_id = 12427 then
	sram_write <= x"02C000C8";
end if;
if first_state_sram_input_id = 12428 then
	sram_write <= x"22EA0220";
end if;
if first_state_sram_input_id = 12429 then
	sram_write <= x"D0ECE000";
end if;
if first_state_sram_input_id = 12430 then
	sram_write <= x"C1040004";
end if;
if first_state_sram_input_id = 12431 then
	sram_write <= x"C1240000";
end if;
if first_state_sram_input_id = 12432 then
	sram_write <= x"C14E0004";
end if;
if first_state_sram_input_id = 12433 then
	sram_write <= x"02800001";
end if;
if first_state_sram_input_id = 12434 then
	sram_write <= x"C45C004C";
end if;
if first_state_sram_input_id = 12435 then
	sram_write <= x"C4DC0050";
end if;
if first_state_sram_input_id = 12436 then
	sram_write <= x"8348C2D4";
end if;
if first_state_sram_input_id = 12437 then
	sram_write <= x"02800002";
end if;
if first_state_sram_input_id = 12438 then
	sram_write <= x"8348C298";
end if;
if first_state_sram_input_id = 12439 then
	sram_write <= x"C51C0054";
end if;
if first_state_sram_input_id = 12440 then
	sram_write <= x"C4BC0058";
end if;
if first_state_sram_input_id = 12441 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12442 then
	sram_write <= x"004E0000";
end if;
if first_state_sram_input_id = 12443 then
	sram_write <= x"00320000";
end if;
if first_state_sram_input_id = 12444 then
	sram_write <= x"03DC0064";
end if;
if first_state_sram_input_id = 12445 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12446 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12447 then
	sram_write <= x"8200400C";
end if;
if first_state_sram_input_id = 12448 then
	sram_write <= x"07DC0064";
end if;
if first_state_sram_input_id = 12449 then
	sram_write <= x"C05C0058";
end if;
if first_state_sram_input_id = 12450 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 12451 then
	sram_write <= x"C09C0054";
end if;
if first_state_sram_input_id = 12452 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 12453 then
	sram_write <= x"8200C2D0";
end if;
if first_state_sram_input_id = 12454 then
	sram_write <= x"C51C0054";
end if;
if first_state_sram_input_id = 12455 then
	sram_write <= x"C4BC0058";
end if;
if first_state_sram_input_id = 12456 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12457 then
	sram_write <= x"004E0000";
end if;
if first_state_sram_input_id = 12458 then
	sram_write <= x"00320000";
end if;
if first_state_sram_input_id = 12459 then
	sram_write <= x"03DC0064";
end if;
if first_state_sram_input_id = 12460 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12461 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12462 then
	sram_write <= x"82003E98";
end if;
if first_state_sram_input_id = 12463 then
	sram_write <= x"07DC0064";
end if;
if first_state_sram_input_id = 12464 then
	sram_write <= x"C05C0058";
end if;
if first_state_sram_input_id = 12465 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 12466 then
	sram_write <= x"C09C0054";
end if;
if first_state_sram_input_id = 12467 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 12468 then
	sram_write <= x"8200C30C";
end if;
if first_state_sram_input_id = 12469 then
	sram_write <= x"C51C0054";
end if;
if first_state_sram_input_id = 12470 then
	sram_write <= x"C4BC0058";
end if;
if first_state_sram_input_id = 12471 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12472 then
	sram_write <= x"004E0000";
end if;
if first_state_sram_input_id = 12473 then
	sram_write <= x"00320000";
end if;
if first_state_sram_input_id = 12474 then
	sram_write <= x"03DC0064";
end if;
if first_state_sram_input_id = 12475 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12476 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12477 then
	sram_write <= x"82003CC4";
end if;
if first_state_sram_input_id = 12478 then
	sram_write <= x"07DC0064";
end if;
if first_state_sram_input_id = 12479 then
	sram_write <= x"C05C0058";
end if;
if first_state_sram_input_id = 12480 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 12481 then
	sram_write <= x"C09C0054";
end if;
if first_state_sram_input_id = 12482 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 12483 then
	sram_write <= x"06240001";
end if;
if first_state_sram_input_id = 12484 then
	sram_write <= x"8620C408";
end if;
if first_state_sram_input_id = 12485 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 12486 then
	sram_write <= x"C07C0050";
end if;
if first_state_sram_input_id = 12487 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 12488 then
	sram_write <= x"C07C004C";
end if;
if first_state_sram_input_id = 12489 then
	sram_write <= x"C0860004";
end if;
if first_state_sram_input_id = 12490 then
	sram_write <= x"C0A60000";
end if;
if first_state_sram_input_id = 12491 then
	sram_write <= x"C0C40004";
end if;
if first_state_sram_input_id = 12492 then
	sram_write <= x"02E00001";
end if;
if first_state_sram_input_id = 12493 then
	sram_write <= x"82CEC3B0";
end if;
if first_state_sram_input_id = 12494 then
	sram_write <= x"02E00002";
end if;
if first_state_sram_input_id = 12495 then
	sram_write <= x"82CEC378";
end if;
if first_state_sram_input_id = 12496 then
	sram_write <= x"C49C005C";
end if;
if first_state_sram_input_id = 12497 then
	sram_write <= x"C43C0060";
end if;
if first_state_sram_input_id = 12498 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12499 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 12500 then
	sram_write <= x"03DC006C";
end if;
if first_state_sram_input_id = 12501 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12502 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12503 then
	sram_write <= x"8200400C";
end if;
if first_state_sram_input_id = 12504 then
	sram_write <= x"07DC006C";
end if;
if first_state_sram_input_id = 12505 then
	sram_write <= x"C05C0060";
end if;
if first_state_sram_input_id = 12506 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 12507 then
	sram_write <= x"C09C005C";
end if;
if first_state_sram_input_id = 12508 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 12509 then
	sram_write <= x"8200C3AC";
end if;
if first_state_sram_input_id = 12510 then
	sram_write <= x"C49C005C";
end if;
if first_state_sram_input_id = 12511 then
	sram_write <= x"C43C0060";
end if;
if first_state_sram_input_id = 12512 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12513 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 12514 then
	sram_write <= x"03DC006C";
end if;
if first_state_sram_input_id = 12515 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12516 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12517 then
	sram_write <= x"82003E98";
end if;
if first_state_sram_input_id = 12518 then
	sram_write <= x"07DC006C";
end if;
if first_state_sram_input_id = 12519 then
	sram_write <= x"C05C0060";
end if;
if first_state_sram_input_id = 12520 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 12521 then
	sram_write <= x"C09C005C";
end if;
if first_state_sram_input_id = 12522 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 12523 then
	sram_write <= x"8200C3E4";
end if;
if first_state_sram_input_id = 12524 then
	sram_write <= x"C49C005C";
end if;
if first_state_sram_input_id = 12525 then
	sram_write <= x"C43C0060";
end if;
if first_state_sram_input_id = 12526 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12527 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 12528 then
	sram_write <= x"03DC006C";
end if;
if first_state_sram_input_id = 12529 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12530 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12531 then
	sram_write <= x"82003CC4";
end if;
if first_state_sram_input_id = 12532 then
	sram_write <= x"07DC006C";
end if;
if first_state_sram_input_id = 12533 then
	sram_write <= x"C05C0060";
end if;
if first_state_sram_input_id = 12534 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 12535 then
	sram_write <= x"C09C005C";
end if;
if first_state_sram_input_id = 12536 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 12537 then
	sram_write <= x"06440001";
end if;
if first_state_sram_input_id = 12538 then
	sram_write <= x"C03C004C";
end if;
if first_state_sram_input_id = 12539 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12540 then
	sram_write <= x"03DC006C";
end if;
if first_state_sram_input_id = 12541 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12542 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12543 then
	sram_write <= x"820042A4";
end if;
if first_state_sram_input_id = 12544 then
	sram_write <= x"07DC006C";
end if;
if first_state_sram_input_id = 12545 then
	sram_write <= x"8200C408";
end if;
if first_state_sram_input_id = 12546 then
	sram_write <= x"8200C40C";
end if;
if first_state_sram_input_id = 12547 then
	sram_write <= x"C03C0048";
end if;
if first_state_sram_input_id = 12548 then
	sram_write <= x"06220001";
end if;
if first_state_sram_input_id = 12549 then
	sram_write <= x"8620C704";
end if;
if first_state_sram_input_id = 12550 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 12551 then
	sram_write <= x"C07C0004";
end if;
if first_state_sram_input_id = 12552 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 12553 then
	sram_write <= x"C09C0000";
end if;
if first_state_sram_input_id = 12554 then
	sram_write <= x"C0880000";
end if;
if first_state_sram_input_id = 12555 then
	sram_write <= x"06880001";
end if;
if first_state_sram_input_id = 12556 then
	sram_write <= x"C43C0064";
end if;
if first_state_sram_input_id = 12557 then
	sram_write <= x"8680C6F4";
end if;
if first_state_sram_input_id = 12558 then
	sram_write <= x"02A000C8";
end if;
if first_state_sram_input_id = 12559 then
	sram_write <= x"22C80220";
end if;
if first_state_sram_input_id = 12560 then
	sram_write <= x"D0CAC000";
end if;
if first_state_sram_input_id = 12561 then
	sram_write <= x"C0E40004";
end if;
if first_state_sram_input_id = 12562 then
	sram_write <= x"C1040000";
end if;
if first_state_sram_input_id = 12563 then
	sram_write <= x"C12C0004";
end if;
if first_state_sram_input_id = 12564 then
	sram_write <= x"03400001";
end if;
if first_state_sram_input_id = 12565 then
	sram_write <= x"C45C0068";
end if;
if first_state_sram_input_id = 12566 then
	sram_write <= x"C4BC006C";
end if;
if first_state_sram_input_id = 12567 then
	sram_write <= x"8334C4E0";
end if;
if first_state_sram_input_id = 12568 then
	sram_write <= x"03400002";
end if;
if first_state_sram_input_id = 12569 then
	sram_write <= x"8334C4A4";
end if;
if first_state_sram_input_id = 12570 then
	sram_write <= x"C4FC0070";
end if;
if first_state_sram_input_id = 12571 then
	sram_write <= x"C49C0074";
end if;
if first_state_sram_input_id = 12572 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12573 then
	sram_write <= x"004C0000";
end if;
if first_state_sram_input_id = 12574 then
	sram_write <= x"00300000";
end if;
if first_state_sram_input_id = 12575 then
	sram_write <= x"03DC0080";
end if;
if first_state_sram_input_id = 12576 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12577 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12578 then
	sram_write <= x"8200400C";
end if;
if first_state_sram_input_id = 12579 then
	sram_write <= x"07DC0080";
end if;
if first_state_sram_input_id = 12580 then
	sram_write <= x"C05C0074";
end if;
if first_state_sram_input_id = 12581 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 12582 then
	sram_write <= x"C09C0070";
end if;
if first_state_sram_input_id = 12583 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 12584 then
	sram_write <= x"8200C4DC";
end if;
if first_state_sram_input_id = 12585 then
	sram_write <= x"C4FC0070";
end if;
if first_state_sram_input_id = 12586 then
	sram_write <= x"C49C0074";
end if;
if first_state_sram_input_id = 12587 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12588 then
	sram_write <= x"004C0000";
end if;
if first_state_sram_input_id = 12589 then
	sram_write <= x"00300000";
end if;
if first_state_sram_input_id = 12590 then
	sram_write <= x"03DC0080";
end if;
if first_state_sram_input_id = 12591 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12592 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12593 then
	sram_write <= x"82003E98";
end if;
if first_state_sram_input_id = 12594 then
	sram_write <= x"07DC0080";
end if;
if first_state_sram_input_id = 12595 then
	sram_write <= x"C05C0074";
end if;
if first_state_sram_input_id = 12596 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 12597 then
	sram_write <= x"C09C0070";
end if;
if first_state_sram_input_id = 12598 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 12599 then
	sram_write <= x"8200C518";
end if;
if first_state_sram_input_id = 12600 then
	sram_write <= x"C4FC0070";
end if;
if first_state_sram_input_id = 12601 then
	sram_write <= x"C49C0074";
end if;
if first_state_sram_input_id = 12602 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12603 then
	sram_write <= x"004C0000";
end if;
if first_state_sram_input_id = 12604 then
	sram_write <= x"00300000";
end if;
if first_state_sram_input_id = 12605 then
	sram_write <= x"03DC0080";
end if;
if first_state_sram_input_id = 12606 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12607 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12608 then
	sram_write <= x"82003CC4";
end if;
if first_state_sram_input_id = 12609 then
	sram_write <= x"07DC0080";
end if;
if first_state_sram_input_id = 12610 then
	sram_write <= x"C05C0074";
end if;
if first_state_sram_input_id = 12611 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 12612 then
	sram_write <= x"C09C0070";
end if;
if first_state_sram_input_id = 12613 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 12614 then
	sram_write <= x"06240001";
end if;
if first_state_sram_input_id = 12615 then
	sram_write <= x"8620C6F0";
end if;
if first_state_sram_input_id = 12616 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 12617 then
	sram_write <= x"C07C006C";
end if;
if first_state_sram_input_id = 12618 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 12619 then
	sram_write <= x"C09C0068";
end if;
if first_state_sram_input_id = 12620 then
	sram_write <= x"C0A80004";
end if;
if first_state_sram_input_id = 12621 then
	sram_write <= x"C0C80000";
end if;
if first_state_sram_input_id = 12622 then
	sram_write <= x"C0E40004";
end if;
if first_state_sram_input_id = 12623 then
	sram_write <= x"03000001";
end if;
if first_state_sram_input_id = 12624 then
	sram_write <= x"82F0C5BC";
end if;
if first_state_sram_input_id = 12625 then
	sram_write <= x"03000002";
end if;
if first_state_sram_input_id = 12626 then
	sram_write <= x"82F0C584";
end if;
if first_state_sram_input_id = 12627 then
	sram_write <= x"C4BC0078";
end if;
if first_state_sram_input_id = 12628 then
	sram_write <= x"C43C007C";
end if;
if first_state_sram_input_id = 12629 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12630 then
	sram_write <= x"002C0000";
end if;
if first_state_sram_input_id = 12631 then
	sram_write <= x"03DC0088";
end if;
if first_state_sram_input_id = 12632 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12633 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12634 then
	sram_write <= x"8200400C";
end if;
if first_state_sram_input_id = 12635 then
	sram_write <= x"07DC0088";
end if;
if first_state_sram_input_id = 12636 then
	sram_write <= x"C05C007C";
end if;
if first_state_sram_input_id = 12637 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 12638 then
	sram_write <= x"C09C0078";
end if;
if first_state_sram_input_id = 12639 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 12640 then
	sram_write <= x"8200C5B8";
end if;
if first_state_sram_input_id = 12641 then
	sram_write <= x"C4BC0078";
end if;
if first_state_sram_input_id = 12642 then
	sram_write <= x"C43C007C";
end if;
if first_state_sram_input_id = 12643 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12644 then
	sram_write <= x"002C0000";
end if;
if first_state_sram_input_id = 12645 then
	sram_write <= x"03DC0088";
end if;
if first_state_sram_input_id = 12646 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12647 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12648 then
	sram_write <= x"82003E98";
end if;
if first_state_sram_input_id = 12649 then
	sram_write <= x"07DC0088";
end if;
if first_state_sram_input_id = 12650 then
	sram_write <= x"C05C007C";
end if;
if first_state_sram_input_id = 12651 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 12652 then
	sram_write <= x"C09C0078";
end if;
if first_state_sram_input_id = 12653 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 12654 then
	sram_write <= x"8200C5F0";
end if;
if first_state_sram_input_id = 12655 then
	sram_write <= x"C4BC0078";
end if;
if first_state_sram_input_id = 12656 then
	sram_write <= x"C43C007C";
end if;
if first_state_sram_input_id = 12657 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12658 then
	sram_write <= x"002C0000";
end if;
if first_state_sram_input_id = 12659 then
	sram_write <= x"03DC0088";
end if;
if first_state_sram_input_id = 12660 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12661 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12662 then
	sram_write <= x"82003CC4";
end if;
if first_state_sram_input_id = 12663 then
	sram_write <= x"07DC0088";
end if;
if first_state_sram_input_id = 12664 then
	sram_write <= x"C05C007C";
end if;
if first_state_sram_input_id = 12665 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 12666 then
	sram_write <= x"C09C0078";
end if;
if first_state_sram_input_id = 12667 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 12668 then
	sram_write <= x"06240001";
end if;
if first_state_sram_input_id = 12669 then
	sram_write <= x"8620C6EC";
end if;
if first_state_sram_input_id = 12670 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 12671 then
	sram_write <= x"C07C006C";
end if;
if first_state_sram_input_id = 12672 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 12673 then
	sram_write <= x"C07C0068";
end if;
if first_state_sram_input_id = 12674 then
	sram_write <= x"C0860004";
end if;
if first_state_sram_input_id = 12675 then
	sram_write <= x"C0A60000";
end if;
if first_state_sram_input_id = 12676 then
	sram_write <= x"C0C40004";
end if;
if first_state_sram_input_id = 12677 then
	sram_write <= x"02E00001";
end if;
if first_state_sram_input_id = 12678 then
	sram_write <= x"82CEC694";
end if;
if first_state_sram_input_id = 12679 then
	sram_write <= x"02E00002";
end if;
if first_state_sram_input_id = 12680 then
	sram_write <= x"82CEC65C";
end if;
if first_state_sram_input_id = 12681 then
	sram_write <= x"C49C0080";
end if;
if first_state_sram_input_id = 12682 then
	sram_write <= x"C43C0084";
end if;
if first_state_sram_input_id = 12683 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12684 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 12685 then
	sram_write <= x"03DC0090";
end if;
if first_state_sram_input_id = 12686 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12687 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12688 then
	sram_write <= x"8200400C";
end if;
if first_state_sram_input_id = 12689 then
	sram_write <= x"07DC0090";
end if;
if first_state_sram_input_id = 12690 then
	sram_write <= x"C05C0084";
end if;
if first_state_sram_input_id = 12691 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 12692 then
	sram_write <= x"C09C0080";
end if;
if first_state_sram_input_id = 12693 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 12694 then
	sram_write <= x"8200C690";
end if;
if first_state_sram_input_id = 12695 then
	sram_write <= x"C49C0080";
end if;
if first_state_sram_input_id = 12696 then
	sram_write <= x"C43C0084";
end if;
if first_state_sram_input_id = 12697 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12698 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 12699 then
	sram_write <= x"03DC0090";
end if;
if first_state_sram_input_id = 12700 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12701 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12702 then
	sram_write <= x"82003E98";
end if;
if first_state_sram_input_id = 12703 then
	sram_write <= x"07DC0090";
end if;
if first_state_sram_input_id = 12704 then
	sram_write <= x"C05C0084";
end if;
if first_state_sram_input_id = 12705 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 12706 then
	sram_write <= x"C09C0080";
end if;
if first_state_sram_input_id = 12707 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 12708 then
	sram_write <= x"8200C6C8";
end if;
if first_state_sram_input_id = 12709 then
	sram_write <= x"C49C0080";
end if;
if first_state_sram_input_id = 12710 then
	sram_write <= x"C43C0084";
end if;
if first_state_sram_input_id = 12711 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12712 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 12713 then
	sram_write <= x"03DC0090";
end if;
if first_state_sram_input_id = 12714 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12715 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12716 then
	sram_write <= x"82003CC4";
end if;
if first_state_sram_input_id = 12717 then
	sram_write <= x"07DC0090";
end if;
if first_state_sram_input_id = 12718 then
	sram_write <= x"C05C0084";
end if;
if first_state_sram_input_id = 12719 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 12720 then
	sram_write <= x"C09C0080";
end if;
if first_state_sram_input_id = 12721 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 12722 then
	sram_write <= x"06440001";
end if;
if first_state_sram_input_id = 12723 then
	sram_write <= x"C03C0068";
end if;
if first_state_sram_input_id = 12724 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12725 then
	sram_write <= x"03DC0090";
end if;
if first_state_sram_input_id = 12726 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12727 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12728 then
	sram_write <= x"820042A4";
end if;
if first_state_sram_input_id = 12729 then
	sram_write <= x"07DC0090";
end if;
if first_state_sram_input_id = 12730 then
	sram_write <= x"8200C6EC";
end if;
if first_state_sram_input_id = 12731 then
	sram_write <= x"8200C6F0";
end if;
if first_state_sram_input_id = 12732 then
	sram_write <= x"8200C6F4";
end if;
if first_state_sram_input_id = 12733 then
	sram_write <= x"C03C0064";
end if;
if first_state_sram_input_id = 12734 then
	sram_write <= x"06420001";
end if;
if first_state_sram_input_id = 12735 then
	sram_write <= x"C03C0004";
end if;
if first_state_sram_input_id = 12736 then
	sram_write <= x"8200BD10";
end if;
if first_state_sram_input_id = 12737 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 12738 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 12739 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 12740 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 12741 then
	sram_write <= x"8620D760";
end if;
if first_state_sram_input_id = 12742 then
	sram_write <= x"02400354";
end if;
if first_state_sram_input_id = 12743 then
	sram_write <= x"22620220";
end if;
if first_state_sram_input_id = 12744 then
	sram_write <= x"D0646000";
end if;
if first_state_sram_input_id = 12745 then
	sram_write <= x"C08601DC";
end if;
if first_state_sram_input_id = 12746 then
	sram_write <= x"02A000C4";
end if;
if first_state_sram_input_id = 12747 then
	sram_write <= x"C0CA0000";
end if;
if first_state_sram_input_id = 12748 then
	sram_write <= x"06CC0001";
end if;
if first_state_sram_input_id = 12749 then
	sram_write <= x"C45C0000";
end if;
if first_state_sram_input_id = 12750 then
	sram_write <= x"C43C0004";
end if;
if first_state_sram_input_id = 12751 then
	sram_write <= x"C4BC0008";
end if;
if first_state_sram_input_id = 12752 then
	sram_write <= x"C47C000C";
end if;
if first_state_sram_input_id = 12753 then
	sram_write <= x"86C0CA04";
end if;
if first_state_sram_input_id = 12754 then
	sram_write <= x"02E000C8";
end if;
if first_state_sram_input_id = 12755 then
	sram_write <= x"230C0220";
end if;
if first_state_sram_input_id = 12756 then
	sram_write <= x"D10F0000";
end if;
if first_state_sram_input_id = 12757 then
	sram_write <= x"C1280004";
end if;
if first_state_sram_input_id = 12758 then
	sram_write <= x"C1480000";
end if;
if first_state_sram_input_id = 12759 then
	sram_write <= x"C0500004";
end if;
if first_state_sram_input_id = 12760 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 12761 then
	sram_write <= x"C49C0010";
end if;
if first_state_sram_input_id = 12762 then
	sram_write <= x"C4FC0014";
end if;
if first_state_sram_input_id = 12763 then
	sram_write <= x"8242C7F0";
end if;
if first_state_sram_input_id = 12764 then
	sram_write <= x"02200002";
end if;
if first_state_sram_input_id = 12765 then
	sram_write <= x"8242C7B4";
end if;
if first_state_sram_input_id = 12766 then
	sram_write <= x"C53C0018";
end if;
if first_state_sram_input_id = 12767 then
	sram_write <= x"C4DC001C";
end if;
if first_state_sram_input_id = 12768 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12769 then
	sram_write <= x"00500000";
end if;
if first_state_sram_input_id = 12770 then
	sram_write <= x"00340000";
end if;
if first_state_sram_input_id = 12771 then
	sram_write <= x"03DC0028";
end if;
if first_state_sram_input_id = 12772 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12773 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12774 then
	sram_write <= x"8200400C";
end if;
if first_state_sram_input_id = 12775 then
	sram_write <= x"07DC0028";
end if;
if first_state_sram_input_id = 12776 then
	sram_write <= x"C05C001C";
end if;
if first_state_sram_input_id = 12777 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 12778 then
	sram_write <= x"C09C0018";
end if;
if first_state_sram_input_id = 12779 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 12780 then
	sram_write <= x"8200C7EC";
end if;
if first_state_sram_input_id = 12781 then
	sram_write <= x"C53C0018";
end if;
if first_state_sram_input_id = 12782 then
	sram_write <= x"C4DC001C";
end if;
if first_state_sram_input_id = 12783 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12784 then
	sram_write <= x"00500000";
end if;
if first_state_sram_input_id = 12785 then
	sram_write <= x"00340000";
end if;
if first_state_sram_input_id = 12786 then
	sram_write <= x"03DC0028";
end if;
if first_state_sram_input_id = 12787 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12788 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12789 then
	sram_write <= x"82003E98";
end if;
if first_state_sram_input_id = 12790 then
	sram_write <= x"07DC0028";
end if;
if first_state_sram_input_id = 12791 then
	sram_write <= x"C05C001C";
end if;
if first_state_sram_input_id = 12792 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 12793 then
	sram_write <= x"C09C0018";
end if;
if first_state_sram_input_id = 12794 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 12795 then
	sram_write <= x"8200C828";
end if;
if first_state_sram_input_id = 12796 then
	sram_write <= x"C53C0018";
end if;
if first_state_sram_input_id = 12797 then
	sram_write <= x"C4DC001C";
end if;
if first_state_sram_input_id = 12798 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12799 then
	sram_write <= x"00500000";
end if;
if first_state_sram_input_id = 12800 then
	sram_write <= x"00340000";
end if;
if first_state_sram_input_id = 12801 then
	sram_write <= x"03DC0028";
end if;
if first_state_sram_input_id = 12802 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12803 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12804 then
	sram_write <= x"82003CC4";
end if;
if first_state_sram_input_id = 12805 then
	sram_write <= x"07DC0028";
end if;
if first_state_sram_input_id = 12806 then
	sram_write <= x"C05C001C";
end if;
if first_state_sram_input_id = 12807 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 12808 then
	sram_write <= x"C09C0018";
end if;
if first_state_sram_input_id = 12809 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 12810 then
	sram_write <= x"06240001";
end if;
if first_state_sram_input_id = 12811 then
	sram_write <= x"8620CA00";
end if;
if first_state_sram_input_id = 12812 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 12813 then
	sram_write <= x"C07C0014";
end if;
if first_state_sram_input_id = 12814 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 12815 then
	sram_write <= x"C09C0010";
end if;
if first_state_sram_input_id = 12816 then
	sram_write <= x"C0A80004";
end if;
if first_state_sram_input_id = 12817 then
	sram_write <= x"C0C80000";
end if;
if first_state_sram_input_id = 12818 then
	sram_write <= x"C0E40004";
end if;
if first_state_sram_input_id = 12819 then
	sram_write <= x"03000001";
end if;
if first_state_sram_input_id = 12820 then
	sram_write <= x"82F0C8CC";
end if;
if first_state_sram_input_id = 12821 then
	sram_write <= x"03000002";
end if;
if first_state_sram_input_id = 12822 then
	sram_write <= x"82F0C894";
end if;
if first_state_sram_input_id = 12823 then
	sram_write <= x"C4BC0020";
end if;
if first_state_sram_input_id = 12824 then
	sram_write <= x"C43C0024";
end if;
if first_state_sram_input_id = 12825 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12826 then
	sram_write <= x"002C0000";
end if;
if first_state_sram_input_id = 12827 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 12828 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12829 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12830 then
	sram_write <= x"8200400C";
end if;
if first_state_sram_input_id = 12831 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 12832 then
	sram_write <= x"C05C0024";
end if;
if first_state_sram_input_id = 12833 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 12834 then
	sram_write <= x"C09C0020";
end if;
if first_state_sram_input_id = 12835 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 12836 then
	sram_write <= x"8200C8C8";
end if;
if first_state_sram_input_id = 12837 then
	sram_write <= x"C4BC0020";
end if;
if first_state_sram_input_id = 12838 then
	sram_write <= x"C43C0024";
end if;
if first_state_sram_input_id = 12839 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12840 then
	sram_write <= x"002C0000";
end if;
if first_state_sram_input_id = 12841 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 12842 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12843 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12844 then
	sram_write <= x"82003E98";
end if;
if first_state_sram_input_id = 12845 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 12846 then
	sram_write <= x"C05C0024";
end if;
if first_state_sram_input_id = 12847 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 12848 then
	sram_write <= x"C09C0020";
end if;
if first_state_sram_input_id = 12849 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 12850 then
	sram_write <= x"8200C900";
end if;
if first_state_sram_input_id = 12851 then
	sram_write <= x"C4BC0020";
end if;
if first_state_sram_input_id = 12852 then
	sram_write <= x"C43C0024";
end if;
if first_state_sram_input_id = 12853 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12854 then
	sram_write <= x"002C0000";
end if;
if first_state_sram_input_id = 12855 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 12856 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12857 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12858 then
	sram_write <= x"82003CC4";
end if;
if first_state_sram_input_id = 12859 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 12860 then
	sram_write <= x"C05C0024";
end if;
if first_state_sram_input_id = 12861 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 12862 then
	sram_write <= x"C09C0020";
end if;
if first_state_sram_input_id = 12863 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 12864 then
	sram_write <= x"06240001";
end if;
if first_state_sram_input_id = 12865 then
	sram_write <= x"8620C9FC";
end if;
if first_state_sram_input_id = 12866 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 12867 then
	sram_write <= x"C07C0014";
end if;
if first_state_sram_input_id = 12868 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 12869 then
	sram_write <= x"C07C0010";
end if;
if first_state_sram_input_id = 12870 then
	sram_write <= x"C0860004";
end if;
if first_state_sram_input_id = 12871 then
	sram_write <= x"C0A60000";
end if;
if first_state_sram_input_id = 12872 then
	sram_write <= x"C0C40004";
end if;
if first_state_sram_input_id = 12873 then
	sram_write <= x"02E00001";
end if;
if first_state_sram_input_id = 12874 then
	sram_write <= x"82CEC9A4";
end if;
if first_state_sram_input_id = 12875 then
	sram_write <= x"02E00002";
end if;
if first_state_sram_input_id = 12876 then
	sram_write <= x"82CEC96C";
end if;
if first_state_sram_input_id = 12877 then
	sram_write <= x"C49C0028";
end if;
if first_state_sram_input_id = 12878 then
	sram_write <= x"C43C002C";
end if;
if first_state_sram_input_id = 12879 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12880 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 12881 then
	sram_write <= x"03DC0038";
end if;
if first_state_sram_input_id = 12882 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12883 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12884 then
	sram_write <= x"8200400C";
end if;
if first_state_sram_input_id = 12885 then
	sram_write <= x"07DC0038";
end if;
if first_state_sram_input_id = 12886 then
	sram_write <= x"C05C002C";
end if;
if first_state_sram_input_id = 12887 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 12888 then
	sram_write <= x"C09C0028";
end if;
if first_state_sram_input_id = 12889 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 12890 then
	sram_write <= x"8200C9A0";
end if;
if first_state_sram_input_id = 12891 then
	sram_write <= x"C49C0028";
end if;
if first_state_sram_input_id = 12892 then
	sram_write <= x"C43C002C";
end if;
if first_state_sram_input_id = 12893 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12894 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 12895 then
	sram_write <= x"03DC0038";
end if;
if first_state_sram_input_id = 12896 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12897 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12898 then
	sram_write <= x"82003E98";
end if;
if first_state_sram_input_id = 12899 then
	sram_write <= x"07DC0038";
end if;
if first_state_sram_input_id = 12900 then
	sram_write <= x"C05C002C";
end if;
if first_state_sram_input_id = 12901 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 12902 then
	sram_write <= x"C09C0028";
end if;
if first_state_sram_input_id = 12903 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 12904 then
	sram_write <= x"8200C9D8";
end if;
if first_state_sram_input_id = 12905 then
	sram_write <= x"C49C0028";
end if;
if first_state_sram_input_id = 12906 then
	sram_write <= x"C43C002C";
end if;
if first_state_sram_input_id = 12907 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12908 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 12909 then
	sram_write <= x"03DC0038";
end if;
if first_state_sram_input_id = 12910 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12911 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12912 then
	sram_write <= x"82003CC4";
end if;
if first_state_sram_input_id = 12913 then
	sram_write <= x"07DC0038";
end if;
if first_state_sram_input_id = 12914 then
	sram_write <= x"C05C002C";
end if;
if first_state_sram_input_id = 12915 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 12916 then
	sram_write <= x"C09C0028";
end if;
if first_state_sram_input_id = 12917 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 12918 then
	sram_write <= x"06440001";
end if;
if first_state_sram_input_id = 12919 then
	sram_write <= x"C03C0010";
end if;
if first_state_sram_input_id = 12920 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12921 then
	sram_write <= x"03DC0038";
end if;
if first_state_sram_input_id = 12922 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12923 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12924 then
	sram_write <= x"820042A4";
end if;
if first_state_sram_input_id = 12925 then
	sram_write <= x"07DC0038";
end if;
if first_state_sram_input_id = 12926 then
	sram_write <= x"8200C9FC";
end if;
if first_state_sram_input_id = 12927 then
	sram_write <= x"8200CA00";
end if;
if first_state_sram_input_id = 12928 then
	sram_write <= x"8200CA04";
end if;
if first_state_sram_input_id = 12929 then
	sram_write <= x"C03C000C";
end if;
if first_state_sram_input_id = 12930 then
	sram_write <= x"C04201D8";
end if;
if first_state_sram_input_id = 12931 then
	sram_write <= x"C07C0008";
end if;
if first_state_sram_input_id = 12932 then
	sram_write <= x"C0860000";
end if;
if first_state_sram_input_id = 12933 then
	sram_write <= x"06880001";
end if;
if first_state_sram_input_id = 12934 then
	sram_write <= x"8680CBFC";
end if;
if first_state_sram_input_id = 12935 then
	sram_write <= x"02A000C8";
end if;
if first_state_sram_input_id = 12936 then
	sram_write <= x"22C80220";
end if;
if first_state_sram_input_id = 12937 then
	sram_write <= x"D0CAC000";
end if;
if first_state_sram_input_id = 12938 then
	sram_write <= x"C0E40004";
end if;
if first_state_sram_input_id = 12939 then
	sram_write <= x"C1040000";
end if;
if first_state_sram_input_id = 12940 then
	sram_write <= x"C12C0004";
end if;
if first_state_sram_input_id = 12941 then
	sram_write <= x"03400001";
end if;
if first_state_sram_input_id = 12942 then
	sram_write <= x"C45C0030";
end if;
if first_state_sram_input_id = 12943 then
	sram_write <= x"C4BC0034";
end if;
if first_state_sram_input_id = 12944 then
	sram_write <= x"8334CAC4";
end if;
if first_state_sram_input_id = 12945 then
	sram_write <= x"03400002";
end if;
if first_state_sram_input_id = 12946 then
	sram_write <= x"8334CA88";
end if;
if first_state_sram_input_id = 12947 then
	sram_write <= x"C4FC0038";
end if;
if first_state_sram_input_id = 12948 then
	sram_write <= x"C49C003C";
end if;
if first_state_sram_input_id = 12949 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12950 then
	sram_write <= x"004C0000";
end if;
if first_state_sram_input_id = 12951 then
	sram_write <= x"00300000";
end if;
if first_state_sram_input_id = 12952 then
	sram_write <= x"03DC0048";
end if;
if first_state_sram_input_id = 12953 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12954 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12955 then
	sram_write <= x"8200400C";
end if;
if first_state_sram_input_id = 12956 then
	sram_write <= x"07DC0048";
end if;
if first_state_sram_input_id = 12957 then
	sram_write <= x"C05C003C";
end if;
if first_state_sram_input_id = 12958 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 12959 then
	sram_write <= x"C09C0038";
end if;
if first_state_sram_input_id = 12960 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 12961 then
	sram_write <= x"8200CAC0";
end if;
if first_state_sram_input_id = 12962 then
	sram_write <= x"C4FC0038";
end if;
if first_state_sram_input_id = 12963 then
	sram_write <= x"C49C003C";
end if;
if first_state_sram_input_id = 12964 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12965 then
	sram_write <= x"004C0000";
end if;
if first_state_sram_input_id = 12966 then
	sram_write <= x"00300000";
end if;
if first_state_sram_input_id = 12967 then
	sram_write <= x"03DC0048";
end if;
if first_state_sram_input_id = 12968 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12969 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12970 then
	sram_write <= x"82003E98";
end if;
if first_state_sram_input_id = 12971 then
	sram_write <= x"07DC0048";
end if;
if first_state_sram_input_id = 12972 then
	sram_write <= x"C05C003C";
end if;
if first_state_sram_input_id = 12973 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 12974 then
	sram_write <= x"C09C0038";
end if;
if first_state_sram_input_id = 12975 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 12976 then
	sram_write <= x"8200CAFC";
end if;
if first_state_sram_input_id = 12977 then
	sram_write <= x"C4FC0038";
end if;
if first_state_sram_input_id = 12978 then
	sram_write <= x"C49C003C";
end if;
if first_state_sram_input_id = 12979 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 12980 then
	sram_write <= x"004C0000";
end if;
if first_state_sram_input_id = 12981 then
	sram_write <= x"00300000";
end if;
if first_state_sram_input_id = 12982 then
	sram_write <= x"03DC0048";
end if;
if first_state_sram_input_id = 12983 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 12984 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 12985 then
	sram_write <= x"82003CC4";
end if;
if first_state_sram_input_id = 12986 then
	sram_write <= x"07DC0048";
end if;
if first_state_sram_input_id = 12987 then
	sram_write <= x"C05C003C";
end if;
if first_state_sram_input_id = 12988 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 12989 then
	sram_write <= x"C09C0038";
end if;
if first_state_sram_input_id = 12990 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 12991 then
	sram_write <= x"06240001";
end if;
if first_state_sram_input_id = 12992 then
	sram_write <= x"8620CBF8";
end if;
if first_state_sram_input_id = 12993 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 12994 then
	sram_write <= x"C07C0034";
end if;
if first_state_sram_input_id = 12995 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 12996 then
	sram_write <= x"C07C0030";
end if;
if first_state_sram_input_id = 12997 then
	sram_write <= x"C0860004";
end if;
if first_state_sram_input_id = 12998 then
	sram_write <= x"C0A60000";
end if;
if first_state_sram_input_id = 12999 then
	sram_write <= x"C0C40004";
end if;
if first_state_sram_input_id = 13000 then
	sram_write <= x"02E00001";
end if;
if first_state_sram_input_id = 13001 then
	sram_write <= x"82CECBA0";
end if;
if first_state_sram_input_id = 13002 then
	sram_write <= x"02E00002";
end if;
if first_state_sram_input_id = 13003 then
	sram_write <= x"82CECB68";
end if;
if first_state_sram_input_id = 13004 then
	sram_write <= x"C49C0040";
end if;
if first_state_sram_input_id = 13005 then
	sram_write <= x"C43C0044";
end if;
if first_state_sram_input_id = 13006 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13007 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 13008 then
	sram_write <= x"03DC0050";
end if;
if first_state_sram_input_id = 13009 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13010 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13011 then
	sram_write <= x"8200400C";
end if;
if first_state_sram_input_id = 13012 then
	sram_write <= x"07DC0050";
end if;
if first_state_sram_input_id = 13013 then
	sram_write <= x"C05C0044";
end if;
if first_state_sram_input_id = 13014 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 13015 then
	sram_write <= x"C09C0040";
end if;
if first_state_sram_input_id = 13016 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 13017 then
	sram_write <= x"8200CB9C";
end if;
if first_state_sram_input_id = 13018 then
	sram_write <= x"C49C0040";
end if;
if first_state_sram_input_id = 13019 then
	sram_write <= x"C43C0044";
end if;
if first_state_sram_input_id = 13020 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13021 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 13022 then
	sram_write <= x"03DC0050";
end if;
if first_state_sram_input_id = 13023 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13024 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13025 then
	sram_write <= x"82003E98";
end if;
if first_state_sram_input_id = 13026 then
	sram_write <= x"07DC0050";
end if;
if first_state_sram_input_id = 13027 then
	sram_write <= x"C05C0044";
end if;
if first_state_sram_input_id = 13028 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 13029 then
	sram_write <= x"C09C0040";
end if;
if first_state_sram_input_id = 13030 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 13031 then
	sram_write <= x"8200CBD4";
end if;
if first_state_sram_input_id = 13032 then
	sram_write <= x"C49C0040";
end if;
if first_state_sram_input_id = 13033 then
	sram_write <= x"C43C0044";
end if;
if first_state_sram_input_id = 13034 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13035 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 13036 then
	sram_write <= x"03DC0050";
end if;
if first_state_sram_input_id = 13037 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13038 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13039 then
	sram_write <= x"82003CC4";
end if;
if first_state_sram_input_id = 13040 then
	sram_write <= x"07DC0050";
end if;
if first_state_sram_input_id = 13041 then
	sram_write <= x"C05C0044";
end if;
if first_state_sram_input_id = 13042 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 13043 then
	sram_write <= x"C09C0040";
end if;
if first_state_sram_input_id = 13044 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 13045 then
	sram_write <= x"06440001";
end if;
if first_state_sram_input_id = 13046 then
	sram_write <= x"C03C0030";
end if;
if first_state_sram_input_id = 13047 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13048 then
	sram_write <= x"03DC0050";
end if;
if first_state_sram_input_id = 13049 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13050 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13051 then
	sram_write <= x"820042A4";
end if;
if first_state_sram_input_id = 13052 then
	sram_write <= x"07DC0050";
end if;
if first_state_sram_input_id = 13053 then
	sram_write <= x"8200CBF8";
end if;
if first_state_sram_input_id = 13054 then
	sram_write <= x"8200CBFC";
end if;
if first_state_sram_input_id = 13055 then
	sram_write <= x"C03C000C";
end if;
if first_state_sram_input_id = 13056 then
	sram_write <= x"C04201D4";
end if;
if first_state_sram_input_id = 13057 then
	sram_write <= x"C07C0008";
end if;
if first_state_sram_input_id = 13058 then
	sram_write <= x"C0860000";
end if;
if first_state_sram_input_id = 13059 then
	sram_write <= x"06880001";
end if;
if first_state_sram_input_id = 13060 then
	sram_write <= x"8680CED0";
end if;
if first_state_sram_input_id = 13061 then
	sram_write <= x"02A000C8";
end if;
if first_state_sram_input_id = 13062 then
	sram_write <= x"22C80220";
end if;
if first_state_sram_input_id = 13063 then
	sram_write <= x"D0CAC000";
end if;
if first_state_sram_input_id = 13064 then
	sram_write <= x"C0E40004";
end if;
if first_state_sram_input_id = 13065 then
	sram_write <= x"C1040000";
end if;
if first_state_sram_input_id = 13066 then
	sram_write <= x"C12C0004";
end if;
if first_state_sram_input_id = 13067 then
	sram_write <= x"03400001";
end if;
if first_state_sram_input_id = 13068 then
	sram_write <= x"C45C0048";
end if;
if first_state_sram_input_id = 13069 then
	sram_write <= x"C4BC004C";
end if;
if first_state_sram_input_id = 13070 then
	sram_write <= x"8334CCBC";
end if;
if first_state_sram_input_id = 13071 then
	sram_write <= x"03400002";
end if;
if first_state_sram_input_id = 13072 then
	sram_write <= x"8334CC80";
end if;
if first_state_sram_input_id = 13073 then
	sram_write <= x"C4FC0050";
end if;
if first_state_sram_input_id = 13074 then
	sram_write <= x"C49C0054";
end if;
if first_state_sram_input_id = 13075 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13076 then
	sram_write <= x"004C0000";
end if;
if first_state_sram_input_id = 13077 then
	sram_write <= x"00300000";
end if;
if first_state_sram_input_id = 13078 then
	sram_write <= x"03DC0060";
end if;
if first_state_sram_input_id = 13079 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13080 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13081 then
	sram_write <= x"8200400C";
end if;
if first_state_sram_input_id = 13082 then
	sram_write <= x"07DC0060";
end if;
if first_state_sram_input_id = 13083 then
	sram_write <= x"C05C0054";
end if;
if first_state_sram_input_id = 13084 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 13085 then
	sram_write <= x"C09C0050";
end if;
if first_state_sram_input_id = 13086 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 13087 then
	sram_write <= x"8200CCB8";
end if;
if first_state_sram_input_id = 13088 then
	sram_write <= x"C4FC0050";
end if;
if first_state_sram_input_id = 13089 then
	sram_write <= x"C49C0054";
end if;
if first_state_sram_input_id = 13090 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13091 then
	sram_write <= x"004C0000";
end if;
if first_state_sram_input_id = 13092 then
	sram_write <= x"00300000";
end if;
if first_state_sram_input_id = 13093 then
	sram_write <= x"03DC0060";
end if;
if first_state_sram_input_id = 13094 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13095 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13096 then
	sram_write <= x"82003E98";
end if;
if first_state_sram_input_id = 13097 then
	sram_write <= x"07DC0060";
end if;
if first_state_sram_input_id = 13098 then
	sram_write <= x"C05C0054";
end if;
if first_state_sram_input_id = 13099 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 13100 then
	sram_write <= x"C09C0050";
end if;
if first_state_sram_input_id = 13101 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 13102 then
	sram_write <= x"8200CCF4";
end if;
if first_state_sram_input_id = 13103 then
	sram_write <= x"C4FC0050";
end if;
if first_state_sram_input_id = 13104 then
	sram_write <= x"C49C0054";
end if;
if first_state_sram_input_id = 13105 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13106 then
	sram_write <= x"004C0000";
end if;
if first_state_sram_input_id = 13107 then
	sram_write <= x"00300000";
end if;
if first_state_sram_input_id = 13108 then
	sram_write <= x"03DC0060";
end if;
if first_state_sram_input_id = 13109 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13110 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13111 then
	sram_write <= x"82003CC4";
end if;
if first_state_sram_input_id = 13112 then
	sram_write <= x"07DC0060";
end if;
if first_state_sram_input_id = 13113 then
	sram_write <= x"C05C0054";
end if;
if first_state_sram_input_id = 13114 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 13115 then
	sram_write <= x"C09C0050";
end if;
if first_state_sram_input_id = 13116 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 13117 then
	sram_write <= x"06240001";
end if;
if first_state_sram_input_id = 13118 then
	sram_write <= x"8620CECC";
end if;
if first_state_sram_input_id = 13119 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 13120 then
	sram_write <= x"C07C004C";
end if;
if first_state_sram_input_id = 13121 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 13122 then
	sram_write <= x"C09C0048";
end if;
if first_state_sram_input_id = 13123 then
	sram_write <= x"C0A80004";
end if;
if first_state_sram_input_id = 13124 then
	sram_write <= x"C0C80000";
end if;
if first_state_sram_input_id = 13125 then
	sram_write <= x"C0E40004";
end if;
if first_state_sram_input_id = 13126 then
	sram_write <= x"03000001";
end if;
if first_state_sram_input_id = 13127 then
	sram_write <= x"82F0CD98";
end if;
if first_state_sram_input_id = 13128 then
	sram_write <= x"03000002";
end if;
if first_state_sram_input_id = 13129 then
	sram_write <= x"82F0CD60";
end if;
if first_state_sram_input_id = 13130 then
	sram_write <= x"C4BC0058";
end if;
if first_state_sram_input_id = 13131 then
	sram_write <= x"C43C005C";
end if;
if first_state_sram_input_id = 13132 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13133 then
	sram_write <= x"002C0000";
end if;
if first_state_sram_input_id = 13134 then
	sram_write <= x"03DC0068";
end if;
if first_state_sram_input_id = 13135 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13136 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13137 then
	sram_write <= x"8200400C";
end if;
if first_state_sram_input_id = 13138 then
	sram_write <= x"07DC0068";
end if;
if first_state_sram_input_id = 13139 then
	sram_write <= x"C05C005C";
end if;
if first_state_sram_input_id = 13140 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 13141 then
	sram_write <= x"C09C0058";
end if;
if first_state_sram_input_id = 13142 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 13143 then
	sram_write <= x"8200CD94";
end if;
if first_state_sram_input_id = 13144 then
	sram_write <= x"C4BC0058";
end if;
if first_state_sram_input_id = 13145 then
	sram_write <= x"C43C005C";
end if;
if first_state_sram_input_id = 13146 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13147 then
	sram_write <= x"002C0000";
end if;
if first_state_sram_input_id = 13148 then
	sram_write <= x"03DC0068";
end if;
if first_state_sram_input_id = 13149 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13150 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13151 then
	sram_write <= x"82003E98";
end if;
if first_state_sram_input_id = 13152 then
	sram_write <= x"07DC0068";
end if;
if first_state_sram_input_id = 13153 then
	sram_write <= x"C05C005C";
end if;
if first_state_sram_input_id = 13154 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 13155 then
	sram_write <= x"C09C0058";
end if;
if first_state_sram_input_id = 13156 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 13157 then
	sram_write <= x"8200CDCC";
end if;
if first_state_sram_input_id = 13158 then
	sram_write <= x"C4BC0058";
end if;
if first_state_sram_input_id = 13159 then
	sram_write <= x"C43C005C";
end if;
if first_state_sram_input_id = 13160 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13161 then
	sram_write <= x"002C0000";
end if;
if first_state_sram_input_id = 13162 then
	sram_write <= x"03DC0068";
end if;
if first_state_sram_input_id = 13163 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13164 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13165 then
	sram_write <= x"82003CC4";
end if;
if first_state_sram_input_id = 13166 then
	sram_write <= x"07DC0068";
end if;
if first_state_sram_input_id = 13167 then
	sram_write <= x"C05C005C";
end if;
if first_state_sram_input_id = 13168 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 13169 then
	sram_write <= x"C09C0058";
end if;
if first_state_sram_input_id = 13170 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 13171 then
	sram_write <= x"06240001";
end if;
if first_state_sram_input_id = 13172 then
	sram_write <= x"8620CEC8";
end if;
if first_state_sram_input_id = 13173 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 13174 then
	sram_write <= x"C07C004C";
end if;
if first_state_sram_input_id = 13175 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 13176 then
	sram_write <= x"C07C0048";
end if;
if first_state_sram_input_id = 13177 then
	sram_write <= x"C0860004";
end if;
if first_state_sram_input_id = 13178 then
	sram_write <= x"C0A60000";
end if;
if first_state_sram_input_id = 13179 then
	sram_write <= x"C0C40004";
end if;
if first_state_sram_input_id = 13180 then
	sram_write <= x"02E00001";
end if;
if first_state_sram_input_id = 13181 then
	sram_write <= x"82CECE70";
end if;
if first_state_sram_input_id = 13182 then
	sram_write <= x"02E00002";
end if;
if first_state_sram_input_id = 13183 then
	sram_write <= x"82CECE38";
end if;
if first_state_sram_input_id = 13184 then
	sram_write <= x"C49C0060";
end if;
if first_state_sram_input_id = 13185 then
	sram_write <= x"C43C0064";
end if;
if first_state_sram_input_id = 13186 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13187 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 13188 then
	sram_write <= x"03DC0070";
end if;
if first_state_sram_input_id = 13189 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13190 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13191 then
	sram_write <= x"8200400C";
end if;
if first_state_sram_input_id = 13192 then
	sram_write <= x"07DC0070";
end if;
if first_state_sram_input_id = 13193 then
	sram_write <= x"C05C0064";
end if;
if first_state_sram_input_id = 13194 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 13195 then
	sram_write <= x"C09C0060";
end if;
if first_state_sram_input_id = 13196 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 13197 then
	sram_write <= x"8200CE6C";
end if;
if first_state_sram_input_id = 13198 then
	sram_write <= x"C49C0060";
end if;
if first_state_sram_input_id = 13199 then
	sram_write <= x"C43C0064";
end if;
if first_state_sram_input_id = 13200 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13201 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 13202 then
	sram_write <= x"03DC0070";
end if;
if first_state_sram_input_id = 13203 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13204 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13205 then
	sram_write <= x"82003E98";
end if;
if first_state_sram_input_id = 13206 then
	sram_write <= x"07DC0070";
end if;
if first_state_sram_input_id = 13207 then
	sram_write <= x"C05C0064";
end if;
if first_state_sram_input_id = 13208 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 13209 then
	sram_write <= x"C09C0060";
end if;
if first_state_sram_input_id = 13210 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 13211 then
	sram_write <= x"8200CEA4";
end if;
if first_state_sram_input_id = 13212 then
	sram_write <= x"C49C0060";
end if;
if first_state_sram_input_id = 13213 then
	sram_write <= x"C43C0064";
end if;
if first_state_sram_input_id = 13214 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13215 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 13216 then
	sram_write <= x"03DC0070";
end if;
if first_state_sram_input_id = 13217 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13218 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13219 then
	sram_write <= x"82003CC4";
end if;
if first_state_sram_input_id = 13220 then
	sram_write <= x"07DC0070";
end if;
if first_state_sram_input_id = 13221 then
	sram_write <= x"C05C0064";
end if;
if first_state_sram_input_id = 13222 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 13223 then
	sram_write <= x"C09C0060";
end if;
if first_state_sram_input_id = 13224 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 13225 then
	sram_write <= x"06440001";
end if;
if first_state_sram_input_id = 13226 then
	sram_write <= x"C03C0048";
end if;
if first_state_sram_input_id = 13227 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13228 then
	sram_write <= x"03DC0070";
end if;
if first_state_sram_input_id = 13229 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13230 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13231 then
	sram_write <= x"820042A4";
end if;
if first_state_sram_input_id = 13232 then
	sram_write <= x"07DC0070";
end if;
if first_state_sram_input_id = 13233 then
	sram_write <= x"8200CEC8";
end if;
if first_state_sram_input_id = 13234 then
	sram_write <= x"8200CECC";
end if;
if first_state_sram_input_id = 13235 then
	sram_write <= x"8200CED0";
end if;
if first_state_sram_input_id = 13236 then
	sram_write <= x"02400074";
end if;
if first_state_sram_input_id = 13237 then
	sram_write <= x"C03C000C";
end if;
if first_state_sram_input_id = 13238 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13239 then
	sram_write <= x"03DC0070";
end if;
if first_state_sram_input_id = 13240 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13241 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13242 then
	sram_write <= x"8200BD10";
end if;
if first_state_sram_input_id = 13243 then
	sram_write <= x"07DC0070";
end if;
if first_state_sram_input_id = 13244 then
	sram_write <= x"C03C0004";
end if;
if first_state_sram_input_id = 13245 then
	sram_write <= x"06220001";
end if;
if first_state_sram_input_id = 13246 then
	sram_write <= x"8620D75C";
end if;
if first_state_sram_input_id = 13247 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 13248 then
	sram_write <= x"C07C0000";
end if;
if first_state_sram_input_id = 13249 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 13250 then
	sram_write <= x"C08401DC";
end if;
if first_state_sram_input_id = 13251 then
	sram_write <= x"C0BC0008";
end if;
if first_state_sram_input_id = 13252 then
	sram_write <= x"C0CA0000";
end if;
if first_state_sram_input_id = 13253 then
	sram_write <= x"06CC0001";
end if;
if first_state_sram_input_id = 13254 then
	sram_write <= x"C43C0068";
end if;
if first_state_sram_input_id = 13255 then
	sram_write <= x"C45C006C";
end if;
if first_state_sram_input_id = 13256 then
	sram_write <= x"86C0D104";
end if;
if first_state_sram_input_id = 13257 then
	sram_write <= x"02E000C8";
end if;
if first_state_sram_input_id = 13258 then
	sram_write <= x"230C0220";
end if;
if first_state_sram_input_id = 13259 then
	sram_write <= x"D10F0000";
end if;
if first_state_sram_input_id = 13260 then
	sram_write <= x"C1280004";
end if;
if first_state_sram_input_id = 13261 then
	sram_write <= x"C1480000";
end if;
if first_state_sram_input_id = 13262 then
	sram_write <= x"C0700004";
end if;
if first_state_sram_input_id = 13263 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 13264 then
	sram_write <= x"C49C0070";
end if;
if first_state_sram_input_id = 13265 then
	sram_write <= x"C4FC0074";
end if;
if first_state_sram_input_id = 13266 then
	sram_write <= x"8262CFCC";
end if;
if first_state_sram_input_id = 13267 then
	sram_write <= x"02200002";
end if;
if first_state_sram_input_id = 13268 then
	sram_write <= x"8262CF90";
end if;
if first_state_sram_input_id = 13269 then
	sram_write <= x"C53C0078";
end if;
if first_state_sram_input_id = 13270 then
	sram_write <= x"C4DC007C";
end if;
if first_state_sram_input_id = 13271 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13272 then
	sram_write <= x"00500000";
end if;
if first_state_sram_input_id = 13273 then
	sram_write <= x"00340000";
end if;
if first_state_sram_input_id = 13274 then
	sram_write <= x"03DC0088";
end if;
if first_state_sram_input_id = 13275 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13276 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13277 then
	sram_write <= x"8200400C";
end if;
if first_state_sram_input_id = 13278 then
	sram_write <= x"07DC0088";
end if;
if first_state_sram_input_id = 13279 then
	sram_write <= x"C05C007C";
end if;
if first_state_sram_input_id = 13280 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 13281 then
	sram_write <= x"C09C0078";
end if;
if first_state_sram_input_id = 13282 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 13283 then
	sram_write <= x"8200CFC8";
end if;
if first_state_sram_input_id = 13284 then
	sram_write <= x"C53C0078";
end if;
if first_state_sram_input_id = 13285 then
	sram_write <= x"C4DC007C";
end if;
if first_state_sram_input_id = 13286 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13287 then
	sram_write <= x"00500000";
end if;
if first_state_sram_input_id = 13288 then
	sram_write <= x"00340000";
end if;
if first_state_sram_input_id = 13289 then
	sram_write <= x"03DC0088";
end if;
if first_state_sram_input_id = 13290 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13291 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13292 then
	sram_write <= x"82003E98";
end if;
if first_state_sram_input_id = 13293 then
	sram_write <= x"07DC0088";
end if;
if first_state_sram_input_id = 13294 then
	sram_write <= x"C05C007C";
end if;
if first_state_sram_input_id = 13295 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 13296 then
	sram_write <= x"C09C0078";
end if;
if first_state_sram_input_id = 13297 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 13298 then
	sram_write <= x"8200D004";
end if;
if first_state_sram_input_id = 13299 then
	sram_write <= x"C53C0078";
end if;
if first_state_sram_input_id = 13300 then
	sram_write <= x"C4DC007C";
end if;
if first_state_sram_input_id = 13301 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13302 then
	sram_write <= x"00500000";
end if;
if first_state_sram_input_id = 13303 then
	sram_write <= x"00340000";
end if;
if first_state_sram_input_id = 13304 then
	sram_write <= x"03DC0088";
end if;
if first_state_sram_input_id = 13305 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13306 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13307 then
	sram_write <= x"82003CC4";
end if;
if first_state_sram_input_id = 13308 then
	sram_write <= x"07DC0088";
end if;
if first_state_sram_input_id = 13309 then
	sram_write <= x"C05C007C";
end if;
if first_state_sram_input_id = 13310 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 13311 then
	sram_write <= x"C09C0078";
end if;
if first_state_sram_input_id = 13312 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 13313 then
	sram_write <= x"06240001";
end if;
if first_state_sram_input_id = 13314 then
	sram_write <= x"8620D100";
end if;
if first_state_sram_input_id = 13315 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 13316 then
	sram_write <= x"C07C0074";
end if;
if first_state_sram_input_id = 13317 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 13318 then
	sram_write <= x"C07C0070";
end if;
if first_state_sram_input_id = 13319 then
	sram_write <= x"C0860004";
end if;
if first_state_sram_input_id = 13320 then
	sram_write <= x"C0A60000";
end if;
if first_state_sram_input_id = 13321 then
	sram_write <= x"C0C40004";
end if;
if first_state_sram_input_id = 13322 then
	sram_write <= x"02E00001";
end if;
if first_state_sram_input_id = 13323 then
	sram_write <= x"82CED0A8";
end if;
if first_state_sram_input_id = 13324 then
	sram_write <= x"02E00002";
end if;
if first_state_sram_input_id = 13325 then
	sram_write <= x"82CED070";
end if;
if first_state_sram_input_id = 13326 then
	sram_write <= x"C49C0080";
end if;
if first_state_sram_input_id = 13327 then
	sram_write <= x"C43C0084";
end if;
if first_state_sram_input_id = 13328 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13329 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 13330 then
	sram_write <= x"03DC0090";
end if;
if first_state_sram_input_id = 13331 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13332 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13333 then
	sram_write <= x"8200400C";
end if;
if first_state_sram_input_id = 13334 then
	sram_write <= x"07DC0090";
end if;
if first_state_sram_input_id = 13335 then
	sram_write <= x"C05C0084";
end if;
if first_state_sram_input_id = 13336 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 13337 then
	sram_write <= x"C09C0080";
end if;
if first_state_sram_input_id = 13338 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 13339 then
	sram_write <= x"8200D0A4";
end if;
if first_state_sram_input_id = 13340 then
	sram_write <= x"C49C0080";
end if;
if first_state_sram_input_id = 13341 then
	sram_write <= x"C43C0084";
end if;
if first_state_sram_input_id = 13342 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13343 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 13344 then
	sram_write <= x"03DC0090";
end if;
if first_state_sram_input_id = 13345 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13346 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13347 then
	sram_write <= x"82003E98";
end if;
if first_state_sram_input_id = 13348 then
	sram_write <= x"07DC0090";
end if;
if first_state_sram_input_id = 13349 then
	sram_write <= x"C05C0084";
end if;
if first_state_sram_input_id = 13350 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 13351 then
	sram_write <= x"C09C0080";
end if;
if first_state_sram_input_id = 13352 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 13353 then
	sram_write <= x"8200D0DC";
end if;
if first_state_sram_input_id = 13354 then
	sram_write <= x"C49C0080";
end if;
if first_state_sram_input_id = 13355 then
	sram_write <= x"C43C0084";
end if;
if first_state_sram_input_id = 13356 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13357 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 13358 then
	sram_write <= x"03DC0090";
end if;
if first_state_sram_input_id = 13359 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13360 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13361 then
	sram_write <= x"82003CC4";
end if;
if first_state_sram_input_id = 13362 then
	sram_write <= x"07DC0090";
end if;
if first_state_sram_input_id = 13363 then
	sram_write <= x"C05C0084";
end if;
if first_state_sram_input_id = 13364 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 13365 then
	sram_write <= x"C09C0080";
end if;
if first_state_sram_input_id = 13366 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 13367 then
	sram_write <= x"06440001";
end if;
if first_state_sram_input_id = 13368 then
	sram_write <= x"C03C0070";
end if;
if first_state_sram_input_id = 13369 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13370 then
	sram_write <= x"03DC0090";
end if;
if first_state_sram_input_id = 13371 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13372 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13373 then
	sram_write <= x"820042A4";
end if;
if first_state_sram_input_id = 13374 then
	sram_write <= x"07DC0090";
end if;
if first_state_sram_input_id = 13375 then
	sram_write <= x"8200D100";
end if;
if first_state_sram_input_id = 13376 then
	sram_write <= x"8200D104";
end if;
if first_state_sram_input_id = 13377 then
	sram_write <= x"C03C006C";
end if;
if first_state_sram_input_id = 13378 then
	sram_write <= x"C04201D8";
end if;
if first_state_sram_input_id = 13379 then
	sram_write <= x"C07C0008";
end if;
if first_state_sram_input_id = 13380 then
	sram_write <= x"C0860000";
end if;
if first_state_sram_input_id = 13381 then
	sram_write <= x"06880001";
end if;
if first_state_sram_input_id = 13382 then
	sram_write <= x"8680D3D8";
end if;
if first_state_sram_input_id = 13383 then
	sram_write <= x"02A000C8";
end if;
if first_state_sram_input_id = 13384 then
	sram_write <= x"22C80220";
end if;
if first_state_sram_input_id = 13385 then
	sram_write <= x"D0CAC000";
end if;
if first_state_sram_input_id = 13386 then
	sram_write <= x"C0E40004";
end if;
if first_state_sram_input_id = 13387 then
	sram_write <= x"C1040000";
end if;
if first_state_sram_input_id = 13388 then
	sram_write <= x"C12C0004";
end if;
if first_state_sram_input_id = 13389 then
	sram_write <= x"03400001";
end if;
if first_state_sram_input_id = 13390 then
	sram_write <= x"C45C0088";
end if;
if first_state_sram_input_id = 13391 then
	sram_write <= x"C4BC008C";
end if;
if first_state_sram_input_id = 13392 then
	sram_write <= x"8334D1C4";
end if;
if first_state_sram_input_id = 13393 then
	sram_write <= x"03400002";
end if;
if first_state_sram_input_id = 13394 then
	sram_write <= x"8334D188";
end if;
if first_state_sram_input_id = 13395 then
	sram_write <= x"C4FC0090";
end if;
if first_state_sram_input_id = 13396 then
	sram_write <= x"C49C0094";
end if;
if first_state_sram_input_id = 13397 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13398 then
	sram_write <= x"004C0000";
end if;
if first_state_sram_input_id = 13399 then
	sram_write <= x"00300000";
end if;
if first_state_sram_input_id = 13400 then
	sram_write <= x"03DC00A0";
end if;
if first_state_sram_input_id = 13401 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13402 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13403 then
	sram_write <= x"8200400C";
end if;
if first_state_sram_input_id = 13404 then
	sram_write <= x"07DC00A0";
end if;
if first_state_sram_input_id = 13405 then
	sram_write <= x"C05C0094";
end if;
if first_state_sram_input_id = 13406 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 13407 then
	sram_write <= x"C09C0090";
end if;
if first_state_sram_input_id = 13408 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 13409 then
	sram_write <= x"8200D1C0";
end if;
if first_state_sram_input_id = 13410 then
	sram_write <= x"C4FC0090";
end if;
if first_state_sram_input_id = 13411 then
	sram_write <= x"C49C0094";
end if;
if first_state_sram_input_id = 13412 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13413 then
	sram_write <= x"004C0000";
end if;
if first_state_sram_input_id = 13414 then
	sram_write <= x"00300000";
end if;
if first_state_sram_input_id = 13415 then
	sram_write <= x"03DC00A0";
end if;
if first_state_sram_input_id = 13416 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13417 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13418 then
	sram_write <= x"82003E98";
end if;
if first_state_sram_input_id = 13419 then
	sram_write <= x"07DC00A0";
end if;
if first_state_sram_input_id = 13420 then
	sram_write <= x"C05C0094";
end if;
if first_state_sram_input_id = 13421 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 13422 then
	sram_write <= x"C09C0090";
end if;
if first_state_sram_input_id = 13423 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 13424 then
	sram_write <= x"8200D1FC";
end if;
if first_state_sram_input_id = 13425 then
	sram_write <= x"C4FC0090";
end if;
if first_state_sram_input_id = 13426 then
	sram_write <= x"C49C0094";
end if;
if first_state_sram_input_id = 13427 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13428 then
	sram_write <= x"004C0000";
end if;
if first_state_sram_input_id = 13429 then
	sram_write <= x"00300000";
end if;
if first_state_sram_input_id = 13430 then
	sram_write <= x"03DC00A0";
end if;
if first_state_sram_input_id = 13431 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13432 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13433 then
	sram_write <= x"82003CC4";
end if;
if first_state_sram_input_id = 13434 then
	sram_write <= x"07DC00A0";
end if;
if first_state_sram_input_id = 13435 then
	sram_write <= x"C05C0094";
end if;
if first_state_sram_input_id = 13436 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 13437 then
	sram_write <= x"C09C0090";
end if;
if first_state_sram_input_id = 13438 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 13439 then
	sram_write <= x"06240001";
end if;
if first_state_sram_input_id = 13440 then
	sram_write <= x"8620D3D4";
end if;
if first_state_sram_input_id = 13441 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 13442 then
	sram_write <= x"C07C008C";
end if;
if first_state_sram_input_id = 13443 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 13444 then
	sram_write <= x"C09C0088";
end if;
if first_state_sram_input_id = 13445 then
	sram_write <= x"C0A80004";
end if;
if first_state_sram_input_id = 13446 then
	sram_write <= x"C0C80000";
end if;
if first_state_sram_input_id = 13447 then
	sram_write <= x"C0E40004";
end if;
if first_state_sram_input_id = 13448 then
	sram_write <= x"03000001";
end if;
if first_state_sram_input_id = 13449 then
	sram_write <= x"82F0D2A0";
end if;
if first_state_sram_input_id = 13450 then
	sram_write <= x"03000002";
end if;
if first_state_sram_input_id = 13451 then
	sram_write <= x"82F0D268";
end if;
if first_state_sram_input_id = 13452 then
	sram_write <= x"C4BC0098";
end if;
if first_state_sram_input_id = 13453 then
	sram_write <= x"C43C009C";
end if;
if first_state_sram_input_id = 13454 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13455 then
	sram_write <= x"002C0000";
end if;
if first_state_sram_input_id = 13456 then
	sram_write <= x"03DC00A8";
end if;
if first_state_sram_input_id = 13457 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13458 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13459 then
	sram_write <= x"8200400C";
end if;
if first_state_sram_input_id = 13460 then
	sram_write <= x"07DC00A8";
end if;
if first_state_sram_input_id = 13461 then
	sram_write <= x"C05C009C";
end if;
if first_state_sram_input_id = 13462 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 13463 then
	sram_write <= x"C09C0098";
end if;
if first_state_sram_input_id = 13464 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 13465 then
	sram_write <= x"8200D29C";
end if;
if first_state_sram_input_id = 13466 then
	sram_write <= x"C4BC0098";
end if;
if first_state_sram_input_id = 13467 then
	sram_write <= x"C43C009C";
end if;
if first_state_sram_input_id = 13468 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13469 then
	sram_write <= x"002C0000";
end if;
if first_state_sram_input_id = 13470 then
	sram_write <= x"03DC00A8";
end if;
if first_state_sram_input_id = 13471 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13472 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13473 then
	sram_write <= x"82003E98";
end if;
if first_state_sram_input_id = 13474 then
	sram_write <= x"07DC00A8";
end if;
if first_state_sram_input_id = 13475 then
	sram_write <= x"C05C009C";
end if;
if first_state_sram_input_id = 13476 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 13477 then
	sram_write <= x"C09C0098";
end if;
if first_state_sram_input_id = 13478 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 13479 then
	sram_write <= x"8200D2D4";
end if;
if first_state_sram_input_id = 13480 then
	sram_write <= x"C4BC0098";
end if;
if first_state_sram_input_id = 13481 then
	sram_write <= x"C43C009C";
end if;
if first_state_sram_input_id = 13482 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13483 then
	sram_write <= x"002C0000";
end if;
if first_state_sram_input_id = 13484 then
	sram_write <= x"03DC00A8";
end if;
if first_state_sram_input_id = 13485 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13486 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13487 then
	sram_write <= x"82003CC4";
end if;
if first_state_sram_input_id = 13488 then
	sram_write <= x"07DC00A8";
end if;
if first_state_sram_input_id = 13489 then
	sram_write <= x"C05C009C";
end if;
if first_state_sram_input_id = 13490 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 13491 then
	sram_write <= x"C09C0098";
end if;
if first_state_sram_input_id = 13492 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 13493 then
	sram_write <= x"06240001";
end if;
if first_state_sram_input_id = 13494 then
	sram_write <= x"8620D3D0";
end if;
if first_state_sram_input_id = 13495 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 13496 then
	sram_write <= x"C07C008C";
end if;
if first_state_sram_input_id = 13497 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 13498 then
	sram_write <= x"C07C0088";
end if;
if first_state_sram_input_id = 13499 then
	sram_write <= x"C0860004";
end if;
if first_state_sram_input_id = 13500 then
	sram_write <= x"C0A60000";
end if;
if first_state_sram_input_id = 13501 then
	sram_write <= x"C0C40004";
end if;
if first_state_sram_input_id = 13502 then
	sram_write <= x"02E00001";
end if;
if first_state_sram_input_id = 13503 then
	sram_write <= x"82CED378";
end if;
if first_state_sram_input_id = 13504 then
	sram_write <= x"02E00002";
end if;
if first_state_sram_input_id = 13505 then
	sram_write <= x"82CED340";
end if;
if first_state_sram_input_id = 13506 then
	sram_write <= x"C49C00A0";
end if;
if first_state_sram_input_id = 13507 then
	sram_write <= x"C43C00A4";
end if;
if first_state_sram_input_id = 13508 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13509 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 13510 then
	sram_write <= x"03DC00B0";
end if;
if first_state_sram_input_id = 13511 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13512 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13513 then
	sram_write <= x"8200400C";
end if;
if first_state_sram_input_id = 13514 then
	sram_write <= x"07DC00B0";
end if;
if first_state_sram_input_id = 13515 then
	sram_write <= x"C05C00A4";
end if;
if first_state_sram_input_id = 13516 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 13517 then
	sram_write <= x"C09C00A0";
end if;
if first_state_sram_input_id = 13518 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 13519 then
	sram_write <= x"8200D374";
end if;
if first_state_sram_input_id = 13520 then
	sram_write <= x"C49C00A0";
end if;
if first_state_sram_input_id = 13521 then
	sram_write <= x"C43C00A4";
end if;
if first_state_sram_input_id = 13522 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13523 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 13524 then
	sram_write <= x"03DC00B0";
end if;
if first_state_sram_input_id = 13525 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13526 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13527 then
	sram_write <= x"82003E98";
end if;
if first_state_sram_input_id = 13528 then
	sram_write <= x"07DC00B0";
end if;
if first_state_sram_input_id = 13529 then
	sram_write <= x"C05C00A4";
end if;
if first_state_sram_input_id = 13530 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 13531 then
	sram_write <= x"C09C00A0";
end if;
if first_state_sram_input_id = 13532 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 13533 then
	sram_write <= x"8200D3AC";
end if;
if first_state_sram_input_id = 13534 then
	sram_write <= x"C49C00A0";
end if;
if first_state_sram_input_id = 13535 then
	sram_write <= x"C43C00A4";
end if;
if first_state_sram_input_id = 13536 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13537 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 13538 then
	sram_write <= x"03DC00B0";
end if;
if first_state_sram_input_id = 13539 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13540 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13541 then
	sram_write <= x"82003CC4";
end if;
if first_state_sram_input_id = 13542 then
	sram_write <= x"07DC00B0";
end if;
if first_state_sram_input_id = 13543 then
	sram_write <= x"C05C00A4";
end if;
if first_state_sram_input_id = 13544 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 13545 then
	sram_write <= x"C09C00A0";
end if;
if first_state_sram_input_id = 13546 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 13547 then
	sram_write <= x"06440001";
end if;
if first_state_sram_input_id = 13548 then
	sram_write <= x"C03C0088";
end if;
if first_state_sram_input_id = 13549 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13550 then
	sram_write <= x"03DC00B0";
end if;
if first_state_sram_input_id = 13551 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13552 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13553 then
	sram_write <= x"820042A4";
end if;
if first_state_sram_input_id = 13554 then
	sram_write <= x"07DC00B0";
end if;
if first_state_sram_input_id = 13555 then
	sram_write <= x"8200D3D0";
end if;
if first_state_sram_input_id = 13556 then
	sram_write <= x"8200D3D4";
end if;
if first_state_sram_input_id = 13557 then
	sram_write <= x"8200D3D8";
end if;
if first_state_sram_input_id = 13558 then
	sram_write <= x"02400075";
end if;
if first_state_sram_input_id = 13559 then
	sram_write <= x"C03C006C";
end if;
if first_state_sram_input_id = 13560 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13561 then
	sram_write <= x"03DC00B0";
end if;
if first_state_sram_input_id = 13562 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13563 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13564 then
	sram_write <= x"8200BD10";
end if;
if first_state_sram_input_id = 13565 then
	sram_write <= x"07DC00B0";
end if;
if first_state_sram_input_id = 13566 then
	sram_write <= x"C03C0068";
end if;
if first_state_sram_input_id = 13567 then
	sram_write <= x"06220001";
end if;
if first_state_sram_input_id = 13568 then
	sram_write <= x"8620D758";
end if;
if first_state_sram_input_id = 13569 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 13570 then
	sram_write <= x"C07C0000";
end if;
if first_state_sram_input_id = 13571 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 13572 then
	sram_write <= x"C08401DC";
end if;
if first_state_sram_input_id = 13573 then
	sram_write <= x"C0BC0008";
end if;
if first_state_sram_input_id = 13574 then
	sram_write <= x"C0AA0000";
end if;
if first_state_sram_input_id = 13575 then
	sram_write <= x"06AA0001";
end if;
if first_state_sram_input_id = 13576 then
	sram_write <= x"C43C00A8";
end if;
if first_state_sram_input_id = 13577 then
	sram_write <= x"C45C00AC";
end if;
if first_state_sram_input_id = 13578 then
	sram_write <= x"86A0D6E8";
end if;
if first_state_sram_input_id = 13579 then
	sram_write <= x"02C000C8";
end if;
if first_state_sram_input_id = 13580 then
	sram_write <= x"22EA0220";
end if;
if first_state_sram_input_id = 13581 then
	sram_write <= x"D0ECE000";
end if;
if first_state_sram_input_id = 13582 then
	sram_write <= x"C1080004";
end if;
if first_state_sram_input_id = 13583 then
	sram_write <= x"C1280000";
end if;
if first_state_sram_input_id = 13584 then
	sram_write <= x"C14E0004";
end if;
if first_state_sram_input_id = 13585 then
	sram_write <= x"02600001";
end if;
if first_state_sram_input_id = 13586 then
	sram_write <= x"C49C00B0";
end if;
if first_state_sram_input_id = 13587 then
	sram_write <= x"C4DC00B4";
end if;
if first_state_sram_input_id = 13588 then
	sram_write <= x"8346D4D4";
end if;
if first_state_sram_input_id = 13589 then
	sram_write <= x"02600002";
end if;
if first_state_sram_input_id = 13590 then
	sram_write <= x"8346D498";
end if;
if first_state_sram_input_id = 13591 then
	sram_write <= x"C51C00B8";
end if;
if first_state_sram_input_id = 13592 then
	sram_write <= x"C4BC00BC";
end if;
if first_state_sram_input_id = 13593 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13594 then
	sram_write <= x"004E0000";
end if;
if first_state_sram_input_id = 13595 then
	sram_write <= x"00320000";
end if;
if first_state_sram_input_id = 13596 then
	sram_write <= x"03DC00C8";
end if;
if first_state_sram_input_id = 13597 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13598 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13599 then
	sram_write <= x"8200400C";
end if;
if first_state_sram_input_id = 13600 then
	sram_write <= x"07DC00C8";
end if;
if first_state_sram_input_id = 13601 then
	sram_write <= x"C05C00BC";
end if;
if first_state_sram_input_id = 13602 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 13603 then
	sram_write <= x"C09C00B8";
end if;
if first_state_sram_input_id = 13604 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 13605 then
	sram_write <= x"8200D4D0";
end if;
if first_state_sram_input_id = 13606 then
	sram_write <= x"C51C00B8";
end if;
if first_state_sram_input_id = 13607 then
	sram_write <= x"C4BC00BC";
end if;
if first_state_sram_input_id = 13608 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13609 then
	sram_write <= x"004E0000";
end if;
if first_state_sram_input_id = 13610 then
	sram_write <= x"00320000";
end if;
if first_state_sram_input_id = 13611 then
	sram_write <= x"03DC00C8";
end if;
if first_state_sram_input_id = 13612 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13613 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13614 then
	sram_write <= x"82003E98";
end if;
if first_state_sram_input_id = 13615 then
	sram_write <= x"07DC00C8";
end if;
if first_state_sram_input_id = 13616 then
	sram_write <= x"C05C00BC";
end if;
if first_state_sram_input_id = 13617 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 13618 then
	sram_write <= x"C09C00B8";
end if;
if first_state_sram_input_id = 13619 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 13620 then
	sram_write <= x"8200D50C";
end if;
if first_state_sram_input_id = 13621 then
	sram_write <= x"C51C00B8";
end if;
if first_state_sram_input_id = 13622 then
	sram_write <= x"C4BC00BC";
end if;
if first_state_sram_input_id = 13623 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13624 then
	sram_write <= x"004E0000";
end if;
if first_state_sram_input_id = 13625 then
	sram_write <= x"00320000";
end if;
if first_state_sram_input_id = 13626 then
	sram_write <= x"03DC00C8";
end if;
if first_state_sram_input_id = 13627 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13628 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13629 then
	sram_write <= x"82003CC4";
end if;
if first_state_sram_input_id = 13630 then
	sram_write <= x"07DC00C8";
end if;
if first_state_sram_input_id = 13631 then
	sram_write <= x"C05C00BC";
end if;
if first_state_sram_input_id = 13632 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 13633 then
	sram_write <= x"C09C00B8";
end if;
if first_state_sram_input_id = 13634 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 13635 then
	sram_write <= x"06240001";
end if;
if first_state_sram_input_id = 13636 then
	sram_write <= x"8620D6E4";
end if;
if first_state_sram_input_id = 13637 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 13638 then
	sram_write <= x"C07C00B4";
end if;
if first_state_sram_input_id = 13639 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 13640 then
	sram_write <= x"C09C00B0";
end if;
if first_state_sram_input_id = 13641 then
	sram_write <= x"C0A80004";
end if;
if first_state_sram_input_id = 13642 then
	sram_write <= x"C0C80000";
end if;
if first_state_sram_input_id = 13643 then
	sram_write <= x"C0E40004";
end if;
if first_state_sram_input_id = 13644 then
	sram_write <= x"03000001";
end if;
if first_state_sram_input_id = 13645 then
	sram_write <= x"82F0D5B0";
end if;
if first_state_sram_input_id = 13646 then
	sram_write <= x"03000002";
end if;
if first_state_sram_input_id = 13647 then
	sram_write <= x"82F0D578";
end if;
if first_state_sram_input_id = 13648 then
	sram_write <= x"C4BC00C0";
end if;
if first_state_sram_input_id = 13649 then
	sram_write <= x"C43C00C4";
end if;
if first_state_sram_input_id = 13650 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13651 then
	sram_write <= x"002C0000";
end if;
if first_state_sram_input_id = 13652 then
	sram_write <= x"03DC00D0";
end if;
if first_state_sram_input_id = 13653 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13654 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13655 then
	sram_write <= x"8200400C";
end if;
if first_state_sram_input_id = 13656 then
	sram_write <= x"07DC00D0";
end if;
if first_state_sram_input_id = 13657 then
	sram_write <= x"C05C00C4";
end if;
if first_state_sram_input_id = 13658 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 13659 then
	sram_write <= x"C09C00C0";
end if;
if first_state_sram_input_id = 13660 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 13661 then
	sram_write <= x"8200D5AC";
end if;
if first_state_sram_input_id = 13662 then
	sram_write <= x"C4BC00C0";
end if;
if first_state_sram_input_id = 13663 then
	sram_write <= x"C43C00C4";
end if;
if first_state_sram_input_id = 13664 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13665 then
	sram_write <= x"002C0000";
end if;
if first_state_sram_input_id = 13666 then
	sram_write <= x"03DC00D0";
end if;
if first_state_sram_input_id = 13667 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13668 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13669 then
	sram_write <= x"82003E98";
end if;
if first_state_sram_input_id = 13670 then
	sram_write <= x"07DC00D0";
end if;
if first_state_sram_input_id = 13671 then
	sram_write <= x"C05C00C4";
end if;
if first_state_sram_input_id = 13672 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 13673 then
	sram_write <= x"C09C00C0";
end if;
if first_state_sram_input_id = 13674 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 13675 then
	sram_write <= x"8200D5E4";
end if;
if first_state_sram_input_id = 13676 then
	sram_write <= x"C4BC00C0";
end if;
if first_state_sram_input_id = 13677 then
	sram_write <= x"C43C00C4";
end if;
if first_state_sram_input_id = 13678 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13679 then
	sram_write <= x"002C0000";
end if;
if first_state_sram_input_id = 13680 then
	sram_write <= x"03DC00D0";
end if;
if first_state_sram_input_id = 13681 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13682 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13683 then
	sram_write <= x"82003CC4";
end if;
if first_state_sram_input_id = 13684 then
	sram_write <= x"07DC00D0";
end if;
if first_state_sram_input_id = 13685 then
	sram_write <= x"C05C00C4";
end if;
if first_state_sram_input_id = 13686 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 13687 then
	sram_write <= x"C09C00C0";
end if;
if first_state_sram_input_id = 13688 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 13689 then
	sram_write <= x"06240001";
end if;
if first_state_sram_input_id = 13690 then
	sram_write <= x"8620D6E0";
end if;
if first_state_sram_input_id = 13691 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 13692 then
	sram_write <= x"C07C00B4";
end if;
if first_state_sram_input_id = 13693 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 13694 then
	sram_write <= x"C07C00B0";
end if;
if first_state_sram_input_id = 13695 then
	sram_write <= x"C0860004";
end if;
if first_state_sram_input_id = 13696 then
	sram_write <= x"C0A60000";
end if;
if first_state_sram_input_id = 13697 then
	sram_write <= x"C0C40004";
end if;
if first_state_sram_input_id = 13698 then
	sram_write <= x"02E00001";
end if;
if first_state_sram_input_id = 13699 then
	sram_write <= x"82CED688";
end if;
if first_state_sram_input_id = 13700 then
	sram_write <= x"02E00002";
end if;
if first_state_sram_input_id = 13701 then
	sram_write <= x"82CED650";
end if;
if first_state_sram_input_id = 13702 then
	sram_write <= x"C49C00C8";
end if;
if first_state_sram_input_id = 13703 then
	sram_write <= x"C43C00CC";
end if;
if first_state_sram_input_id = 13704 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13705 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 13706 then
	sram_write <= x"03DC00D8";
end if;
if first_state_sram_input_id = 13707 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13708 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13709 then
	sram_write <= x"8200400C";
end if;
if first_state_sram_input_id = 13710 then
	sram_write <= x"07DC00D8";
end if;
if first_state_sram_input_id = 13711 then
	sram_write <= x"C05C00CC";
end if;
if first_state_sram_input_id = 13712 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 13713 then
	sram_write <= x"C09C00C8";
end if;
if first_state_sram_input_id = 13714 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 13715 then
	sram_write <= x"8200D684";
end if;
if first_state_sram_input_id = 13716 then
	sram_write <= x"C49C00C8";
end if;
if first_state_sram_input_id = 13717 then
	sram_write <= x"C43C00CC";
end if;
if first_state_sram_input_id = 13718 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13719 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 13720 then
	sram_write <= x"03DC00D8";
end if;
if first_state_sram_input_id = 13721 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13722 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13723 then
	sram_write <= x"82003E98";
end if;
if first_state_sram_input_id = 13724 then
	sram_write <= x"07DC00D8";
end if;
if first_state_sram_input_id = 13725 then
	sram_write <= x"C05C00CC";
end if;
if first_state_sram_input_id = 13726 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 13727 then
	sram_write <= x"C09C00C8";
end if;
if first_state_sram_input_id = 13728 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 13729 then
	sram_write <= x"8200D6BC";
end if;
if first_state_sram_input_id = 13730 then
	sram_write <= x"C49C00C8";
end if;
if first_state_sram_input_id = 13731 then
	sram_write <= x"C43C00CC";
end if;
if first_state_sram_input_id = 13732 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13733 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 13734 then
	sram_write <= x"03DC00D8";
end if;
if first_state_sram_input_id = 13735 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13736 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13737 then
	sram_write <= x"82003CC4";
end if;
if first_state_sram_input_id = 13738 then
	sram_write <= x"07DC00D8";
end if;
if first_state_sram_input_id = 13739 then
	sram_write <= x"C05C00CC";
end if;
if first_state_sram_input_id = 13740 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 13741 then
	sram_write <= x"C09C00C8";
end if;
if first_state_sram_input_id = 13742 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 13743 then
	sram_write <= x"06440001";
end if;
if first_state_sram_input_id = 13744 then
	sram_write <= x"C03C00B0";
end if;
if first_state_sram_input_id = 13745 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13746 then
	sram_write <= x"03DC00D8";
end if;
if first_state_sram_input_id = 13747 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13748 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13749 then
	sram_write <= x"820042A4";
end if;
if first_state_sram_input_id = 13750 then
	sram_write <= x"07DC00D8";
end if;
if first_state_sram_input_id = 13751 then
	sram_write <= x"8200D6E0";
end if;
if first_state_sram_input_id = 13752 then
	sram_write <= x"8200D6E4";
end if;
if first_state_sram_input_id = 13753 then
	sram_write <= x"8200D6E8";
end if;
if first_state_sram_input_id = 13754 then
	sram_write <= x"02400076";
end if;
if first_state_sram_input_id = 13755 then
	sram_write <= x"C03C00AC";
end if;
if first_state_sram_input_id = 13756 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13757 then
	sram_write <= x"03DC00D8";
end if;
if first_state_sram_input_id = 13758 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13759 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13760 then
	sram_write <= x"8200BD10";
end if;
if first_state_sram_input_id = 13761 then
	sram_write <= x"07DC00D8";
end if;
if first_state_sram_input_id = 13762 then
	sram_write <= x"C03C00A8";
end if;
if first_state_sram_input_id = 13763 then
	sram_write <= x"06220001";
end if;
if first_state_sram_input_id = 13764 then
	sram_write <= x"8620D754";
end if;
if first_state_sram_input_id = 13765 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 13766 then
	sram_write <= x"C07C0000";
end if;
if first_state_sram_input_id = 13767 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 13768 then
	sram_write <= x"02600077";
end if;
if first_state_sram_input_id = 13769 then
	sram_write <= x"C43C00D0";
end if;
if first_state_sram_input_id = 13770 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13771 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 13772 then
	sram_write <= x"00460000";
end if;
if first_state_sram_input_id = 13773 then
	sram_write <= x"03DC00DC";
end if;
if first_state_sram_input_id = 13774 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13775 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13776 then
	sram_write <= x"8200BD10";
end if;
if first_state_sram_input_id = 13777 then
	sram_write <= x"07DC00DC";
end if;
if first_state_sram_input_id = 13778 then
	sram_write <= x"C03C00D0";
end if;
if first_state_sram_input_id = 13779 then
	sram_write <= x"06220001";
end if;
if first_state_sram_input_id = 13780 then
	sram_write <= x"8200C714";
end if;
if first_state_sram_input_id = 13781 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 13782 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 13783 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 13784 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 13785 then
	sram_write <= x"22220220";
end if;
if first_state_sram_input_id = 13786 then
	sram_write <= x"02600640";
end if;
if first_state_sram_input_id = 13787 then
	sram_write <= x"C0860000";
end if;
if first_state_sram_input_id = 13788 then
	sram_write <= x"C82000A8";
end if;
if first_state_sram_input_id = 13789 then
	sram_write <= x"C044001C";
end if;
if first_state_sram_input_id = 13790 then
	sram_write <= x"C8440000";
end if;
if first_state_sram_input_id = 13791 then
	sram_write <= x"44224000";
end if;
if first_state_sram_input_id = 13792 then
	sram_write <= x"024001D0";
end if;
if first_state_sram_input_id = 13793 then
	sram_write <= x"C8440000";
end if;
if first_state_sram_input_id = 13794 then
	sram_write <= x"44404000";
end if;
if first_state_sram_input_id = 13795 then
	sram_write <= x"C8640004";
end if;
if first_state_sram_input_id = 13796 then
	sram_write <= x"44606000";
end if;
if first_state_sram_input_id = 13797 then
	sram_write <= x"C8840008";
end if;
if first_state_sram_input_id = 13798 then
	sram_write <= x"44808000";
end if;
if first_state_sram_input_id = 13799 then
	sram_write <= x"02A20001";
end if;
if first_state_sram_input_id = 13800 then
	sram_write <= x"C8A40000";
end if;
if first_state_sram_input_id = 13801 then
	sram_write <= x"02C00003";
end if;
if first_state_sram_input_id = 13802 then
	sram_write <= x"40C00000";
end if;
if first_state_sram_input_id = 13803 then
	sram_write <= x"C47C0000";
end if;
if first_state_sram_input_id = 13804 then
	sram_write <= x"CC5C0008";
end if;
if first_state_sram_input_id = 13805 then
	sram_write <= x"CCDC0010";
end if;
if first_state_sram_input_id = 13806 then
	sram_write <= x"C45C0018";
end if;
if first_state_sram_input_id = 13807 then
	sram_write <= x"C43C001C";
end if;
if first_state_sram_input_id = 13808 then
	sram_write <= x"C49C0020";
end if;
if first_state_sram_input_id = 13809 then
	sram_write <= x"C4BC0024";
end if;
if first_state_sram_input_id = 13810 then
	sram_write <= x"CC3C0028";
end if;
if first_state_sram_input_id = 13811 then
	sram_write <= x"CC9C0030";
end if;
if first_state_sram_input_id = 13812 then
	sram_write <= x"CC7C0038";
end if;
if first_state_sram_input_id = 13813 then
	sram_write <= x"CCBC0040";
end if;
if first_state_sram_input_id = 13814 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13815 then
	sram_write <= x"002C0000";
end if;
if first_state_sram_input_id = 13816 then
	sram_write <= x"4020C000";
end if;
if first_state_sram_input_id = 13817 then
	sram_write <= x"03DC0050";
end if;
if first_state_sram_input_id = 13818 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13819 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13820 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 13821 then
	sram_write <= x"07DC0050";
end if;
if first_state_sram_input_id = 13822 then
	sram_write <= x"00420000";
end if;
if first_state_sram_input_id = 13823 then
	sram_write <= x"022000C4";
end if;
if first_state_sram_input_id = 13824 then
	sram_write <= x"C0620000";
end if;
if first_state_sram_input_id = 13825 then
	sram_write <= x"C43C0048";
end if;
if first_state_sram_input_id = 13826 then
	sram_write <= x"C45C004C";
end if;
if first_state_sram_input_id = 13827 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13828 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 13829 then
	sram_write <= x"03DC0058";
end if;
if first_state_sram_input_id = 13830 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13831 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13832 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 13833 then
	sram_write <= x"07DC0058";
end if;
if first_state_sram_input_id = 13834 then
	sram_write <= x"005A0000";
end if;
if first_state_sram_input_id = 13835 then
	sram_write <= x"03BA0008";
end if;
if first_state_sram_input_id = 13836 then
	sram_write <= x"C4240004";
end if;
if first_state_sram_input_id = 13837 then
	sram_write <= x"C07C004C";
end if;
if first_state_sram_input_id = 13838 then
	sram_write <= x"C4640000";
end if;
if first_state_sram_input_id = 13839 then
	sram_write <= x"C83C0040";
end if;
if first_state_sram_input_id = 13840 then
	sram_write <= x"CC260000";
end if;
if first_state_sram_input_id = 13841 then
	sram_write <= x"C83C0038";
end if;
if first_state_sram_input_id = 13842 then
	sram_write <= x"CC260004";
end if;
if first_state_sram_input_id = 13843 then
	sram_write <= x"C85C0030";
end if;
if first_state_sram_input_id = 13844 then
	sram_write <= x"CC460008";
end if;
if first_state_sram_input_id = 13845 then
	sram_write <= x"C09C0048";
end if;
if first_state_sram_input_id = 13846 then
	sram_write <= x"C0A80000";
end if;
if first_state_sram_input_id = 13847 then
	sram_write <= x"06AA0001";
end if;
if first_state_sram_input_id = 13848 then
	sram_write <= x"C45C0050";
end if;
if first_state_sram_input_id = 13849 then
	sram_write <= x"86A0DB00";
end if;
if first_state_sram_input_id = 13850 then
	sram_write <= x"02C000C8";
end if;
if first_state_sram_input_id = 13851 then
	sram_write <= x"22EA0220";
end if;
if first_state_sram_input_id = 13852 then
	sram_write <= x"D0ECE000";
end if;
if first_state_sram_input_id = 13853 then
	sram_write <= x"C10E0004";
end if;
if first_state_sram_input_id = 13854 then
	sram_write <= x"03200001";
end if;
if first_state_sram_input_id = 13855 then
	sram_write <= x"C4DC0054";
end if;
if first_state_sram_input_id = 13856 then
	sram_write <= x"8312D904";
end if;
if first_state_sram_input_id = 13857 then
	sram_write <= x"03200002";
end if;
if first_state_sram_input_id = 13858 then
	sram_write <= x"8312D8C8";
end if;
if first_state_sram_input_id = 13859 then
	sram_write <= x"C43C0058";
end if;
if first_state_sram_input_id = 13860 then
	sram_write <= x"C4BC005C";
end if;
if first_state_sram_input_id = 13861 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13862 then
	sram_write <= x"004E0000";
end if;
if first_state_sram_input_id = 13863 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 13864 then
	sram_write <= x"03DC0068";
end if;
if first_state_sram_input_id = 13865 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13866 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13867 then
	sram_write <= x"8200400C";
end if;
if first_state_sram_input_id = 13868 then
	sram_write <= x"07DC0068";
end if;
if first_state_sram_input_id = 13869 then
	sram_write <= x"C05C005C";
end if;
if first_state_sram_input_id = 13870 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 13871 then
	sram_write <= x"C09C0058";
end if;
if first_state_sram_input_id = 13872 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 13873 then
	sram_write <= x"8200D900";
end if;
if first_state_sram_input_id = 13874 then
	sram_write <= x"C43C0058";
end if;
if first_state_sram_input_id = 13875 then
	sram_write <= x"C4BC005C";
end if;
if first_state_sram_input_id = 13876 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13877 then
	sram_write <= x"004E0000";
end if;
if first_state_sram_input_id = 13878 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 13879 then
	sram_write <= x"03DC0068";
end if;
if first_state_sram_input_id = 13880 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13881 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13882 then
	sram_write <= x"82003E98";
end if;
if first_state_sram_input_id = 13883 then
	sram_write <= x"07DC0068";
end if;
if first_state_sram_input_id = 13884 then
	sram_write <= x"C05C005C";
end if;
if first_state_sram_input_id = 13885 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 13886 then
	sram_write <= x"C09C0058";
end if;
if first_state_sram_input_id = 13887 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 13888 then
	sram_write <= x"8200D93C";
end if;
if first_state_sram_input_id = 13889 then
	sram_write <= x"C43C0058";
end if;
if first_state_sram_input_id = 13890 then
	sram_write <= x"C4BC005C";
end if;
if first_state_sram_input_id = 13891 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13892 then
	sram_write <= x"004E0000";
end if;
if first_state_sram_input_id = 13893 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 13894 then
	sram_write <= x"03DC0068";
end if;
if first_state_sram_input_id = 13895 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13896 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13897 then
	sram_write <= x"82003CC4";
end if;
if first_state_sram_input_id = 13898 then
	sram_write <= x"07DC0068";
end if;
if first_state_sram_input_id = 13899 then
	sram_write <= x"C05C005C";
end if;
if first_state_sram_input_id = 13900 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 13901 then
	sram_write <= x"C09C0058";
end if;
if first_state_sram_input_id = 13902 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 13903 then
	sram_write <= x"06240001";
end if;
if first_state_sram_input_id = 13904 then
	sram_write <= x"8620DAFC";
end if;
if first_state_sram_input_id = 13905 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 13906 then
	sram_write <= x"C07C0054";
end if;
if first_state_sram_input_id = 13907 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 13908 then
	sram_write <= x"C0A40004";
end if;
if first_state_sram_input_id = 13909 then
	sram_write <= x"02C00001";
end if;
if first_state_sram_input_id = 13910 then
	sram_write <= x"82ACD9D4";
end if;
if first_state_sram_input_id = 13911 then
	sram_write <= x"02C00002";
end if;
if first_state_sram_input_id = 13912 then
	sram_write <= x"82ACD99C";
end if;
if first_state_sram_input_id = 13913 then
	sram_write <= x"C0BC004C";
end if;
if first_state_sram_input_id = 13914 then
	sram_write <= x"C43C0060";
end if;
if first_state_sram_input_id = 13915 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13916 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 13917 then
	sram_write <= x"03DC006C";
end if;
if first_state_sram_input_id = 13918 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13919 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13920 then
	sram_write <= x"8200400C";
end if;
if first_state_sram_input_id = 13921 then
	sram_write <= x"07DC006C";
end if;
if first_state_sram_input_id = 13922 then
	sram_write <= x"C05C0060";
end if;
if first_state_sram_input_id = 13923 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 13924 then
	sram_write <= x"C09C0058";
end if;
if first_state_sram_input_id = 13925 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 13926 then
	sram_write <= x"8200D9D0";
end if;
if first_state_sram_input_id = 13927 then
	sram_write <= x"C0BC004C";
end if;
if first_state_sram_input_id = 13928 then
	sram_write <= x"C43C0060";
end if;
if first_state_sram_input_id = 13929 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13930 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 13931 then
	sram_write <= x"03DC006C";
end if;
if first_state_sram_input_id = 13932 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13933 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13934 then
	sram_write <= x"82003E98";
end if;
if first_state_sram_input_id = 13935 then
	sram_write <= x"07DC006C";
end if;
if first_state_sram_input_id = 13936 then
	sram_write <= x"C05C0060";
end if;
if first_state_sram_input_id = 13937 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 13938 then
	sram_write <= x"C09C0058";
end if;
if first_state_sram_input_id = 13939 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 13940 then
	sram_write <= x"8200DA08";
end if;
if first_state_sram_input_id = 13941 then
	sram_write <= x"C0BC004C";
end if;
if first_state_sram_input_id = 13942 then
	sram_write <= x"C43C0060";
end if;
if first_state_sram_input_id = 13943 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13944 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 13945 then
	sram_write <= x"03DC006C";
end if;
if first_state_sram_input_id = 13946 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13947 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13948 then
	sram_write <= x"82003CC4";
end if;
if first_state_sram_input_id = 13949 then
	sram_write <= x"07DC006C";
end if;
if first_state_sram_input_id = 13950 then
	sram_write <= x"C05C0060";
end if;
if first_state_sram_input_id = 13951 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 13952 then
	sram_write <= x"C09C0058";
end if;
if first_state_sram_input_id = 13953 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 13954 then
	sram_write <= x"06240001";
end if;
if first_state_sram_input_id = 13955 then
	sram_write <= x"8620DAF8";
end if;
if first_state_sram_input_id = 13956 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 13957 then
	sram_write <= x"C07C0054";
end if;
if first_state_sram_input_id = 13958 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 13959 then
	sram_write <= x"C0640004";
end if;
if first_state_sram_input_id = 13960 then
	sram_write <= x"02A00001";
end if;
if first_state_sram_input_id = 13961 then
	sram_write <= x"826ADAA0";
end if;
if first_state_sram_input_id = 13962 then
	sram_write <= x"02A00002";
end if;
if first_state_sram_input_id = 13963 then
	sram_write <= x"826ADA68";
end if;
if first_state_sram_input_id = 13964 then
	sram_write <= x"C07C004C";
end if;
if first_state_sram_input_id = 13965 then
	sram_write <= x"C43C0064";
end if;
if first_state_sram_input_id = 13966 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13967 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 13968 then
	sram_write <= x"03DC0070";
end if;
if first_state_sram_input_id = 13969 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13970 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13971 then
	sram_write <= x"8200400C";
end if;
if first_state_sram_input_id = 13972 then
	sram_write <= x"07DC0070";
end if;
if first_state_sram_input_id = 13973 then
	sram_write <= x"C05C0064";
end if;
if first_state_sram_input_id = 13974 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 13975 then
	sram_write <= x"C09C0058";
end if;
if first_state_sram_input_id = 13976 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 13977 then
	sram_write <= x"8200DA9C";
end if;
if first_state_sram_input_id = 13978 then
	sram_write <= x"C07C004C";
end if;
if first_state_sram_input_id = 13979 then
	sram_write <= x"C43C0064";
end if;
if first_state_sram_input_id = 13980 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13981 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 13982 then
	sram_write <= x"03DC0070";
end if;
if first_state_sram_input_id = 13983 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13984 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13985 then
	sram_write <= x"82003E98";
end if;
if first_state_sram_input_id = 13986 then
	sram_write <= x"07DC0070";
end if;
if first_state_sram_input_id = 13987 then
	sram_write <= x"C05C0064";
end if;
if first_state_sram_input_id = 13988 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 13989 then
	sram_write <= x"C09C0058";
end if;
if first_state_sram_input_id = 13990 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 13991 then
	sram_write <= x"8200DAD4";
end if;
if first_state_sram_input_id = 13992 then
	sram_write <= x"C07C004C";
end if;
if first_state_sram_input_id = 13993 then
	sram_write <= x"C43C0064";
end if;
if first_state_sram_input_id = 13994 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 13995 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 13996 then
	sram_write <= x"03DC0070";
end if;
if first_state_sram_input_id = 13997 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 13998 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 13999 then
	sram_write <= x"82003CC4";
end if;
if first_state_sram_input_id = 14000 then
	sram_write <= x"07DC0070";
end if;
if first_state_sram_input_id = 14001 then
	sram_write <= x"C05C0064";
end if;
if first_state_sram_input_id = 14002 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 14003 then
	sram_write <= x"C09C0058";
end if;
if first_state_sram_input_id = 14004 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 14005 then
	sram_write <= x"06440001";
end if;
if first_state_sram_input_id = 14006 then
	sram_write <= x"C03C0050";
end if;
if first_state_sram_input_id = 14007 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14008 then
	sram_write <= x"03DC0070";
end if;
if first_state_sram_input_id = 14009 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14010 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14011 then
	sram_write <= x"820042A4";
end if;
if first_state_sram_input_id = 14012 then
	sram_write <= x"07DC0070";
end if;
if first_state_sram_input_id = 14013 then
	sram_write <= x"8200DAF8";
end if;
if first_state_sram_input_id = 14014 then
	sram_write <= x"8200DAFC";
end if;
if first_state_sram_input_id = 14015 then
	sram_write <= x"8200DB00";
end if;
if first_state_sram_input_id = 14016 then
	sram_write <= x"02200370";
end if;
if first_state_sram_input_id = 14017 then
	sram_write <= x"005A0000";
end if;
if first_state_sram_input_id = 14018 then
	sram_write <= x"03BA000C";
end if;
if first_state_sram_input_id = 14019 then
	sram_write <= x"C83C0028";
end if;
if first_state_sram_input_id = 14020 then
	sram_write <= x"CC240008";
end if;
if first_state_sram_input_id = 14021 then
	sram_write <= x"C07C0050";
end if;
if first_state_sram_input_id = 14022 then
	sram_write <= x"C4640004";
end if;
if first_state_sram_input_id = 14023 then
	sram_write <= x"C07C0024";
end if;
if first_state_sram_input_id = 14024 then
	sram_write <= x"C4640000";
end if;
if first_state_sram_input_id = 14025 then
	sram_write <= x"C07C0020";
end if;
if first_state_sram_input_id = 14026 then
	sram_write <= x"22860220";
end if;
if first_state_sram_input_id = 14027 then
	sram_write <= x"D4428000";
end if;
if first_state_sram_input_id = 14028 then
	sram_write <= x"02460001";
end if;
if first_state_sram_input_id = 14029 then
	sram_write <= x"C09C001C";
end if;
if first_state_sram_input_id = 14030 then
	sram_write <= x"02A80002";
end if;
if first_state_sram_input_id = 14031 then
	sram_write <= x"C0DC0018";
end if;
if first_state_sram_input_id = 14032 then
	sram_write <= x"C84C0004";
end if;
if first_state_sram_input_id = 14033 then
	sram_write <= x"02E00003";
end if;
if first_state_sram_input_id = 14034 then
	sram_write <= x"C87C0010";
end if;
if first_state_sram_input_id = 14035 then
	sram_write <= x"C43C0068";
end if;
if first_state_sram_input_id = 14036 then
	sram_write <= x"C45C006C";
end if;
if first_state_sram_input_id = 14037 then
	sram_write <= x"C4BC0070";
end if;
if first_state_sram_input_id = 14038 then
	sram_write <= x"CC5C0078";
end if;
if first_state_sram_input_id = 14039 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14040 then
	sram_write <= x"002E0000";
end if;
if first_state_sram_input_id = 14041 then
	sram_write <= x"40206000";
end if;
if first_state_sram_input_id = 14042 then
	sram_write <= x"03DC0088";
end if;
if first_state_sram_input_id = 14043 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14044 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14045 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 14046 then
	sram_write <= x"07DC0088";
end if;
if first_state_sram_input_id = 14047 then
	sram_write <= x"00420000";
end if;
if first_state_sram_input_id = 14048 then
	sram_write <= x"C03C0048";
end if;
if first_state_sram_input_id = 14049 then
	sram_write <= x"C0620000";
end if;
if first_state_sram_input_id = 14050 then
	sram_write <= x"C45C0080";
end if;
if first_state_sram_input_id = 14051 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14052 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 14053 then
	sram_write <= x"03DC008C";
end if;
if first_state_sram_input_id = 14054 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14055 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14056 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 14057 then
	sram_write <= x"07DC008C";
end if;
if first_state_sram_input_id = 14058 then
	sram_write <= x"005A0000";
end if;
if first_state_sram_input_id = 14059 then
	sram_write <= x"03BA0008";
end if;
if first_state_sram_input_id = 14060 then
	sram_write <= x"C4240004";
end if;
if first_state_sram_input_id = 14061 then
	sram_write <= x"C07C0080";
end if;
if first_state_sram_input_id = 14062 then
	sram_write <= x"C4640000";
end if;
if first_state_sram_input_id = 14063 then
	sram_write <= x"C83C0008";
end if;
if first_state_sram_input_id = 14064 then
	sram_write <= x"CC260000";
end if;
if first_state_sram_input_id = 14065 then
	sram_write <= x"C85C0078";
end if;
if first_state_sram_input_id = 14066 then
	sram_write <= x"CC460004";
end if;
if first_state_sram_input_id = 14067 then
	sram_write <= x"C85C0030";
end if;
if first_state_sram_input_id = 14068 then
	sram_write <= x"CC460008";
end if;
if first_state_sram_input_id = 14069 then
	sram_write <= x"C09C0048";
end if;
if first_state_sram_input_id = 14070 then
	sram_write <= x"C0A80000";
end if;
if first_state_sram_input_id = 14071 then
	sram_write <= x"06AA0001";
end if;
if first_state_sram_input_id = 14072 then
	sram_write <= x"C45C0084";
end if;
if first_state_sram_input_id = 14073 then
	sram_write <= x"86A0DE80";
end if;
if first_state_sram_input_id = 14074 then
	sram_write <= x"02C000C8";
end if;
if first_state_sram_input_id = 14075 then
	sram_write <= x"22EA0220";
end if;
if first_state_sram_input_id = 14076 then
	sram_write <= x"D0ECE000";
end if;
if first_state_sram_input_id = 14077 then
	sram_write <= x"C10E0004";
end if;
if first_state_sram_input_id = 14078 then
	sram_write <= x"03200001";
end if;
if first_state_sram_input_id = 14079 then
	sram_write <= x"C4DC0088";
end if;
if first_state_sram_input_id = 14080 then
	sram_write <= x"8312DC84";
end if;
if first_state_sram_input_id = 14081 then
	sram_write <= x"03200002";
end if;
if first_state_sram_input_id = 14082 then
	sram_write <= x"8312DC48";
end if;
if first_state_sram_input_id = 14083 then
	sram_write <= x"C43C008C";
end if;
if first_state_sram_input_id = 14084 then
	sram_write <= x"C4BC0090";
end if;
if first_state_sram_input_id = 14085 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14086 then
	sram_write <= x"004E0000";
end if;
if first_state_sram_input_id = 14087 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 14088 then
	sram_write <= x"03DC009C";
end if;
if first_state_sram_input_id = 14089 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14090 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14091 then
	sram_write <= x"8200400C";
end if;
if first_state_sram_input_id = 14092 then
	sram_write <= x"07DC009C";
end if;
if first_state_sram_input_id = 14093 then
	sram_write <= x"C05C0090";
end if;
if first_state_sram_input_id = 14094 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 14095 then
	sram_write <= x"C09C008C";
end if;
if first_state_sram_input_id = 14096 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 14097 then
	sram_write <= x"8200DC80";
end if;
if first_state_sram_input_id = 14098 then
	sram_write <= x"C43C008C";
end if;
if first_state_sram_input_id = 14099 then
	sram_write <= x"C4BC0090";
end if;
if first_state_sram_input_id = 14100 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14101 then
	sram_write <= x"004E0000";
end if;
if first_state_sram_input_id = 14102 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 14103 then
	sram_write <= x"03DC009C";
end if;
if first_state_sram_input_id = 14104 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14105 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14106 then
	sram_write <= x"82003E98";
end if;
if first_state_sram_input_id = 14107 then
	sram_write <= x"07DC009C";
end if;
if first_state_sram_input_id = 14108 then
	sram_write <= x"C05C0090";
end if;
if first_state_sram_input_id = 14109 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 14110 then
	sram_write <= x"C09C008C";
end if;
if first_state_sram_input_id = 14111 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 14112 then
	sram_write <= x"8200DCBC";
end if;
if first_state_sram_input_id = 14113 then
	sram_write <= x"C43C008C";
end if;
if first_state_sram_input_id = 14114 then
	sram_write <= x"C4BC0090";
end if;
if first_state_sram_input_id = 14115 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14116 then
	sram_write <= x"004E0000";
end if;
if first_state_sram_input_id = 14117 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 14118 then
	sram_write <= x"03DC009C";
end if;
if first_state_sram_input_id = 14119 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14120 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14121 then
	sram_write <= x"82003CC4";
end if;
if first_state_sram_input_id = 14122 then
	sram_write <= x"07DC009C";
end if;
if first_state_sram_input_id = 14123 then
	sram_write <= x"C05C0090";
end if;
if first_state_sram_input_id = 14124 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 14125 then
	sram_write <= x"C09C008C";
end if;
if first_state_sram_input_id = 14126 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 14127 then
	sram_write <= x"06240001";
end if;
if first_state_sram_input_id = 14128 then
	sram_write <= x"8620DE7C";
end if;
if first_state_sram_input_id = 14129 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 14130 then
	sram_write <= x"C07C0088";
end if;
if first_state_sram_input_id = 14131 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 14132 then
	sram_write <= x"C0A40004";
end if;
if first_state_sram_input_id = 14133 then
	sram_write <= x"02C00001";
end if;
if first_state_sram_input_id = 14134 then
	sram_write <= x"82ACDD54";
end if;
if first_state_sram_input_id = 14135 then
	sram_write <= x"02C00002";
end if;
if first_state_sram_input_id = 14136 then
	sram_write <= x"82ACDD1C";
end if;
if first_state_sram_input_id = 14137 then
	sram_write <= x"C0BC0080";
end if;
if first_state_sram_input_id = 14138 then
	sram_write <= x"C43C0094";
end if;
if first_state_sram_input_id = 14139 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14140 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 14141 then
	sram_write <= x"03DC00A0";
end if;
if first_state_sram_input_id = 14142 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14143 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14144 then
	sram_write <= x"8200400C";
end if;
if first_state_sram_input_id = 14145 then
	sram_write <= x"07DC00A0";
end if;
if first_state_sram_input_id = 14146 then
	sram_write <= x"C05C0094";
end if;
if first_state_sram_input_id = 14147 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 14148 then
	sram_write <= x"C09C008C";
end if;
if first_state_sram_input_id = 14149 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 14150 then
	sram_write <= x"8200DD50";
end if;
if first_state_sram_input_id = 14151 then
	sram_write <= x"C0BC0080";
end if;
if first_state_sram_input_id = 14152 then
	sram_write <= x"C43C0094";
end if;
if first_state_sram_input_id = 14153 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14154 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 14155 then
	sram_write <= x"03DC00A0";
end if;
if first_state_sram_input_id = 14156 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14157 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14158 then
	sram_write <= x"82003E98";
end if;
if first_state_sram_input_id = 14159 then
	sram_write <= x"07DC00A0";
end if;
if first_state_sram_input_id = 14160 then
	sram_write <= x"C05C0094";
end if;
if first_state_sram_input_id = 14161 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 14162 then
	sram_write <= x"C09C008C";
end if;
if first_state_sram_input_id = 14163 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 14164 then
	sram_write <= x"8200DD88";
end if;
if first_state_sram_input_id = 14165 then
	sram_write <= x"C0BC0080";
end if;
if first_state_sram_input_id = 14166 then
	sram_write <= x"C43C0094";
end if;
if first_state_sram_input_id = 14167 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14168 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 14169 then
	sram_write <= x"03DC00A0";
end if;
if first_state_sram_input_id = 14170 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14171 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14172 then
	sram_write <= x"82003CC4";
end if;
if first_state_sram_input_id = 14173 then
	sram_write <= x"07DC00A0";
end if;
if first_state_sram_input_id = 14174 then
	sram_write <= x"C05C0094";
end if;
if first_state_sram_input_id = 14175 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 14176 then
	sram_write <= x"C09C008C";
end if;
if first_state_sram_input_id = 14177 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 14178 then
	sram_write <= x"06240001";
end if;
if first_state_sram_input_id = 14179 then
	sram_write <= x"8620DE78";
end if;
if first_state_sram_input_id = 14180 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 14181 then
	sram_write <= x"C07C0088";
end if;
if first_state_sram_input_id = 14182 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 14183 then
	sram_write <= x"C0640004";
end if;
if first_state_sram_input_id = 14184 then
	sram_write <= x"02A00001";
end if;
if first_state_sram_input_id = 14185 then
	sram_write <= x"826ADE20";
end if;
if first_state_sram_input_id = 14186 then
	sram_write <= x"02A00002";
end if;
if first_state_sram_input_id = 14187 then
	sram_write <= x"826ADDE8";
end if;
if first_state_sram_input_id = 14188 then
	sram_write <= x"C07C0080";
end if;
if first_state_sram_input_id = 14189 then
	sram_write <= x"C43C0098";
end if;
if first_state_sram_input_id = 14190 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14191 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 14192 then
	sram_write <= x"03DC00A4";
end if;
if first_state_sram_input_id = 14193 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14194 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14195 then
	sram_write <= x"8200400C";
end if;
if first_state_sram_input_id = 14196 then
	sram_write <= x"07DC00A4";
end if;
if first_state_sram_input_id = 14197 then
	sram_write <= x"C05C0098";
end if;
if first_state_sram_input_id = 14198 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 14199 then
	sram_write <= x"C09C008C";
end if;
if first_state_sram_input_id = 14200 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 14201 then
	sram_write <= x"8200DE1C";
end if;
if first_state_sram_input_id = 14202 then
	sram_write <= x"C07C0080";
end if;
if first_state_sram_input_id = 14203 then
	sram_write <= x"C43C0098";
end if;
if first_state_sram_input_id = 14204 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14205 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 14206 then
	sram_write <= x"03DC00A4";
end if;
if first_state_sram_input_id = 14207 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14208 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14209 then
	sram_write <= x"82003E98";
end if;
if first_state_sram_input_id = 14210 then
	sram_write <= x"07DC00A4";
end if;
if first_state_sram_input_id = 14211 then
	sram_write <= x"C05C0098";
end if;
if first_state_sram_input_id = 14212 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 14213 then
	sram_write <= x"C09C008C";
end if;
if first_state_sram_input_id = 14214 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 14215 then
	sram_write <= x"8200DE54";
end if;
if first_state_sram_input_id = 14216 then
	sram_write <= x"C07C0080";
end if;
if first_state_sram_input_id = 14217 then
	sram_write <= x"C43C0098";
end if;
if first_state_sram_input_id = 14218 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14219 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 14220 then
	sram_write <= x"03DC00A4";
end if;
if first_state_sram_input_id = 14221 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14222 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14223 then
	sram_write <= x"82003CC4";
end if;
if first_state_sram_input_id = 14224 then
	sram_write <= x"07DC00A4";
end if;
if first_state_sram_input_id = 14225 then
	sram_write <= x"C05C0098";
end if;
if first_state_sram_input_id = 14226 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 14227 then
	sram_write <= x"C09C008C";
end if;
if first_state_sram_input_id = 14228 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 14229 then
	sram_write <= x"06440001";
end if;
if first_state_sram_input_id = 14230 then
	sram_write <= x"C03C0084";
end if;
if first_state_sram_input_id = 14231 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14232 then
	sram_write <= x"03DC00A4";
end if;
if first_state_sram_input_id = 14233 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14234 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14235 then
	sram_write <= x"820042A4";
end if;
if first_state_sram_input_id = 14236 then
	sram_write <= x"07DC00A4";
end if;
if first_state_sram_input_id = 14237 then
	sram_write <= x"8200DE78";
end if;
if first_state_sram_input_id = 14238 then
	sram_write <= x"8200DE7C";
end if;
if first_state_sram_input_id = 14239 then
	sram_write <= x"8200DE80";
end if;
if first_state_sram_input_id = 14240 then
	sram_write <= x"003A0000";
end if;
if first_state_sram_input_id = 14241 then
	sram_write <= x"03BA000C";
end if;
if first_state_sram_input_id = 14242 then
	sram_write <= x"C83C0028";
end if;
if first_state_sram_input_id = 14243 then
	sram_write <= x"CC220008";
end if;
if first_state_sram_input_id = 14244 then
	sram_write <= x"C05C0084";
end if;
if first_state_sram_input_id = 14245 then
	sram_write <= x"C4420004";
end if;
if first_state_sram_input_id = 14246 then
	sram_write <= x"C05C0070";
end if;
if first_state_sram_input_id = 14247 then
	sram_write <= x"C4420000";
end if;
if first_state_sram_input_id = 14248 then
	sram_write <= x"C05C006C";
end if;
if first_state_sram_input_id = 14249 then
	sram_write <= x"22440220";
end if;
if first_state_sram_input_id = 14250 then
	sram_write <= x"C07C0068";
end if;
if first_state_sram_input_id = 14251 then
	sram_write <= x"D4264000";
end if;
if first_state_sram_input_id = 14252 then
	sram_write <= x"C03C0020";
end if;
if first_state_sram_input_id = 14253 then
	sram_write <= x"02420002";
end if;
if first_state_sram_input_id = 14254 then
	sram_write <= x"C09C001C";
end if;
if first_state_sram_input_id = 14255 then
	sram_write <= x"02880003";
end if;
if first_state_sram_input_id = 14256 then
	sram_write <= x"C0BC0018";
end if;
if first_state_sram_input_id = 14257 then
	sram_write <= x"C84A0008";
end if;
if first_state_sram_input_id = 14258 then
	sram_write <= x"02A00003";
end if;
if first_state_sram_input_id = 14259 then
	sram_write <= x"C87C0010";
end if;
if first_state_sram_input_id = 14260 then
	sram_write <= x"C45C009C";
end if;
if first_state_sram_input_id = 14261 then
	sram_write <= x"C49C00A0";
end if;
if first_state_sram_input_id = 14262 then
	sram_write <= x"CC5C00A8";
end if;
if first_state_sram_input_id = 14263 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14264 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 14265 then
	sram_write <= x"40206000";
end if;
if first_state_sram_input_id = 14266 then
	sram_write <= x"03DC00B8";
end if;
if first_state_sram_input_id = 14267 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14268 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14269 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 14270 then
	sram_write <= x"07DC00B8";
end if;
if first_state_sram_input_id = 14271 then
	sram_write <= x"00420000";
end if;
if first_state_sram_input_id = 14272 then
	sram_write <= x"C03C0048";
end if;
if first_state_sram_input_id = 14273 then
	sram_write <= x"C0620000";
end if;
if first_state_sram_input_id = 14274 then
	sram_write <= x"C45C00B0";
end if;
if first_state_sram_input_id = 14275 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14276 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 14277 then
	sram_write <= x"03DC00BC";
end if;
if first_state_sram_input_id = 14278 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14279 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14280 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 14281 then
	sram_write <= x"07DC00BC";
end if;
if first_state_sram_input_id = 14282 then
	sram_write <= x"005A0000";
end if;
if first_state_sram_input_id = 14283 then
	sram_write <= x"03BA0008";
end if;
if first_state_sram_input_id = 14284 then
	sram_write <= x"C4240004";
end if;
if first_state_sram_input_id = 14285 then
	sram_write <= x"C07C00B0";
end if;
if first_state_sram_input_id = 14286 then
	sram_write <= x"C4640000";
end if;
if first_state_sram_input_id = 14287 then
	sram_write <= x"C83C0008";
end if;
if first_state_sram_input_id = 14288 then
	sram_write <= x"CC260000";
end if;
if first_state_sram_input_id = 14289 then
	sram_write <= x"C83C0038";
end if;
if first_state_sram_input_id = 14290 then
	sram_write <= x"CC260004";
end if;
if first_state_sram_input_id = 14291 then
	sram_write <= x"C83C00A8";
end if;
if first_state_sram_input_id = 14292 then
	sram_write <= x"CC260008";
end if;
if first_state_sram_input_id = 14293 then
	sram_write <= x"C09C0048";
end if;
if first_state_sram_input_id = 14294 then
	sram_write <= x"C0880000";
end if;
if first_state_sram_input_id = 14295 then
	sram_write <= x"06880001";
end if;
if first_state_sram_input_id = 14296 then
	sram_write <= x"C45C00B4";
end if;
if first_state_sram_input_id = 14297 then
	sram_write <= x"8680E200";
end if;
if first_state_sram_input_id = 14298 then
	sram_write <= x"02A000C8";
end if;
if first_state_sram_input_id = 14299 then
	sram_write <= x"22C80220";
end if;
if first_state_sram_input_id = 14300 then
	sram_write <= x"D0CAC000";
end if;
if first_state_sram_input_id = 14301 then
	sram_write <= x"C0EC0004";
end if;
if first_state_sram_input_id = 14302 then
	sram_write <= x"03000001";
end if;
if first_state_sram_input_id = 14303 then
	sram_write <= x"C4BC00B8";
end if;
if first_state_sram_input_id = 14304 then
	sram_write <= x"82F0E004";
end if;
if first_state_sram_input_id = 14305 then
	sram_write <= x"03000002";
end if;
if first_state_sram_input_id = 14306 then
	sram_write <= x"82F0DFC8";
end if;
if first_state_sram_input_id = 14307 then
	sram_write <= x"C43C00BC";
end if;
if first_state_sram_input_id = 14308 then
	sram_write <= x"C49C00C0";
end if;
if first_state_sram_input_id = 14309 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14310 then
	sram_write <= x"004C0000";
end if;
if first_state_sram_input_id = 14311 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 14312 then
	sram_write <= x"03DC00CC";
end if;
if first_state_sram_input_id = 14313 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14314 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14315 then
	sram_write <= x"8200400C";
end if;
if first_state_sram_input_id = 14316 then
	sram_write <= x"07DC00CC";
end if;
if first_state_sram_input_id = 14317 then
	sram_write <= x"C05C00C0";
end if;
if first_state_sram_input_id = 14318 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 14319 then
	sram_write <= x"C09C00BC";
end if;
if first_state_sram_input_id = 14320 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 14321 then
	sram_write <= x"8200E000";
end if;
if first_state_sram_input_id = 14322 then
	sram_write <= x"C43C00BC";
end if;
if first_state_sram_input_id = 14323 then
	sram_write <= x"C49C00C0";
end if;
if first_state_sram_input_id = 14324 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14325 then
	sram_write <= x"004C0000";
end if;
if first_state_sram_input_id = 14326 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 14327 then
	sram_write <= x"03DC00CC";
end if;
if first_state_sram_input_id = 14328 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14329 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14330 then
	sram_write <= x"82003E98";
end if;
if first_state_sram_input_id = 14331 then
	sram_write <= x"07DC00CC";
end if;
if first_state_sram_input_id = 14332 then
	sram_write <= x"C05C00C0";
end if;
if first_state_sram_input_id = 14333 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 14334 then
	sram_write <= x"C09C00BC";
end if;
if first_state_sram_input_id = 14335 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 14336 then
	sram_write <= x"8200E03C";
end if;
if first_state_sram_input_id = 14337 then
	sram_write <= x"C43C00BC";
end if;
if first_state_sram_input_id = 14338 then
	sram_write <= x"C49C00C0";
end if;
if first_state_sram_input_id = 14339 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14340 then
	sram_write <= x"004C0000";
end if;
if first_state_sram_input_id = 14341 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 14342 then
	sram_write <= x"03DC00CC";
end if;
if first_state_sram_input_id = 14343 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14344 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14345 then
	sram_write <= x"82003CC4";
end if;
if first_state_sram_input_id = 14346 then
	sram_write <= x"07DC00CC";
end if;
if first_state_sram_input_id = 14347 then
	sram_write <= x"C05C00C0";
end if;
if first_state_sram_input_id = 14348 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 14349 then
	sram_write <= x"C09C00BC";
end if;
if first_state_sram_input_id = 14350 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 14351 then
	sram_write <= x"06240001";
end if;
if first_state_sram_input_id = 14352 then
	sram_write <= x"8620E1FC";
end if;
if first_state_sram_input_id = 14353 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 14354 then
	sram_write <= x"C07C00B8";
end if;
if first_state_sram_input_id = 14355 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 14356 then
	sram_write <= x"C0A40004";
end if;
if first_state_sram_input_id = 14357 then
	sram_write <= x"02C00001";
end if;
if first_state_sram_input_id = 14358 then
	sram_write <= x"82ACE0D4";
end if;
if first_state_sram_input_id = 14359 then
	sram_write <= x"02C00002";
end if;
if first_state_sram_input_id = 14360 then
	sram_write <= x"82ACE09C";
end if;
if first_state_sram_input_id = 14361 then
	sram_write <= x"C0BC00B0";
end if;
if first_state_sram_input_id = 14362 then
	sram_write <= x"C43C00C4";
end if;
if first_state_sram_input_id = 14363 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14364 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 14365 then
	sram_write <= x"03DC00D0";
end if;
if first_state_sram_input_id = 14366 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14367 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14368 then
	sram_write <= x"8200400C";
end if;
if first_state_sram_input_id = 14369 then
	sram_write <= x"07DC00D0";
end if;
if first_state_sram_input_id = 14370 then
	sram_write <= x"C05C00C4";
end if;
if first_state_sram_input_id = 14371 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 14372 then
	sram_write <= x"C09C00BC";
end if;
if first_state_sram_input_id = 14373 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 14374 then
	sram_write <= x"8200E0D0";
end if;
if first_state_sram_input_id = 14375 then
	sram_write <= x"C0BC00B0";
end if;
if first_state_sram_input_id = 14376 then
	sram_write <= x"C43C00C4";
end if;
if first_state_sram_input_id = 14377 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14378 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 14379 then
	sram_write <= x"03DC00D0";
end if;
if first_state_sram_input_id = 14380 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14381 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14382 then
	sram_write <= x"82003E98";
end if;
if first_state_sram_input_id = 14383 then
	sram_write <= x"07DC00D0";
end if;
if first_state_sram_input_id = 14384 then
	sram_write <= x"C05C00C4";
end if;
if first_state_sram_input_id = 14385 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 14386 then
	sram_write <= x"C09C00BC";
end if;
if first_state_sram_input_id = 14387 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 14388 then
	sram_write <= x"8200E108";
end if;
if first_state_sram_input_id = 14389 then
	sram_write <= x"C0BC00B0";
end if;
if first_state_sram_input_id = 14390 then
	sram_write <= x"C43C00C4";
end if;
if first_state_sram_input_id = 14391 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14392 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 14393 then
	sram_write <= x"03DC00D0";
end if;
if first_state_sram_input_id = 14394 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14395 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14396 then
	sram_write <= x"82003CC4";
end if;
if first_state_sram_input_id = 14397 then
	sram_write <= x"07DC00D0";
end if;
if first_state_sram_input_id = 14398 then
	sram_write <= x"C05C00C4";
end if;
if first_state_sram_input_id = 14399 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 14400 then
	sram_write <= x"C09C00BC";
end if;
if first_state_sram_input_id = 14401 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 14402 then
	sram_write <= x"06240001";
end if;
if first_state_sram_input_id = 14403 then
	sram_write <= x"8620E1F8";
end if;
if first_state_sram_input_id = 14404 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 14405 then
	sram_write <= x"C07C00B8";
end if;
if first_state_sram_input_id = 14406 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 14407 then
	sram_write <= x"C0640004";
end if;
if first_state_sram_input_id = 14408 then
	sram_write <= x"02A00001";
end if;
if first_state_sram_input_id = 14409 then
	sram_write <= x"826AE1A0";
end if;
if first_state_sram_input_id = 14410 then
	sram_write <= x"02A00002";
end if;
if first_state_sram_input_id = 14411 then
	sram_write <= x"826AE168";
end if;
if first_state_sram_input_id = 14412 then
	sram_write <= x"C07C00B0";
end if;
if first_state_sram_input_id = 14413 then
	sram_write <= x"C43C00C8";
end if;
if first_state_sram_input_id = 14414 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14415 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 14416 then
	sram_write <= x"03DC00D4";
end if;
if first_state_sram_input_id = 14417 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14418 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14419 then
	sram_write <= x"8200400C";
end if;
if first_state_sram_input_id = 14420 then
	sram_write <= x"07DC00D4";
end if;
if first_state_sram_input_id = 14421 then
	sram_write <= x"C05C00C8";
end if;
if first_state_sram_input_id = 14422 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 14423 then
	sram_write <= x"C09C00BC";
end if;
if first_state_sram_input_id = 14424 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 14425 then
	sram_write <= x"8200E19C";
end if;
if first_state_sram_input_id = 14426 then
	sram_write <= x"C07C00B0";
end if;
if first_state_sram_input_id = 14427 then
	sram_write <= x"C43C00C8";
end if;
if first_state_sram_input_id = 14428 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14429 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 14430 then
	sram_write <= x"03DC00D4";
end if;
if first_state_sram_input_id = 14431 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14432 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14433 then
	sram_write <= x"82003E98";
end if;
if first_state_sram_input_id = 14434 then
	sram_write <= x"07DC00D4";
end if;
if first_state_sram_input_id = 14435 then
	sram_write <= x"C05C00C8";
end if;
if first_state_sram_input_id = 14436 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 14437 then
	sram_write <= x"C09C00BC";
end if;
if first_state_sram_input_id = 14438 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 14439 then
	sram_write <= x"8200E1D4";
end if;
if first_state_sram_input_id = 14440 then
	sram_write <= x"C07C00B0";
end if;
if first_state_sram_input_id = 14441 then
	sram_write <= x"C43C00C8";
end if;
if first_state_sram_input_id = 14442 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14443 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 14444 then
	sram_write <= x"03DC00D4";
end if;
if first_state_sram_input_id = 14445 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14446 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14447 then
	sram_write <= x"82003CC4";
end if;
if first_state_sram_input_id = 14448 then
	sram_write <= x"07DC00D4";
end if;
if first_state_sram_input_id = 14449 then
	sram_write <= x"C05C00C8";
end if;
if first_state_sram_input_id = 14450 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 14451 then
	sram_write <= x"C09C00BC";
end if;
if first_state_sram_input_id = 14452 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 14453 then
	sram_write <= x"06440001";
end if;
if first_state_sram_input_id = 14454 then
	sram_write <= x"C03C00B4";
end if;
if first_state_sram_input_id = 14455 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14456 then
	sram_write <= x"03DC00D4";
end if;
if first_state_sram_input_id = 14457 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14458 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14459 then
	sram_write <= x"820042A4";
end if;
if first_state_sram_input_id = 14460 then
	sram_write <= x"07DC00D4";
end if;
if first_state_sram_input_id = 14461 then
	sram_write <= x"8200E1F8";
end if;
if first_state_sram_input_id = 14462 then
	sram_write <= x"8200E1FC";
end if;
if first_state_sram_input_id = 14463 then
	sram_write <= x"8200E200";
end if;
if first_state_sram_input_id = 14464 then
	sram_write <= x"003A0000";
end if;
if first_state_sram_input_id = 14465 then
	sram_write <= x"03BA000C";
end if;
if first_state_sram_input_id = 14466 then
	sram_write <= x"C83C0028";
end if;
if first_state_sram_input_id = 14467 then
	sram_write <= x"CC220008";
end if;
if first_state_sram_input_id = 14468 then
	sram_write <= x"C05C00B4";
end if;
if first_state_sram_input_id = 14469 then
	sram_write <= x"C4420004";
end if;
if first_state_sram_input_id = 14470 then
	sram_write <= x"C05C00A0";
end if;
if first_state_sram_input_id = 14471 then
	sram_write <= x"C4420000";
end if;
if first_state_sram_input_id = 14472 then
	sram_write <= x"C05C009C";
end if;
if first_state_sram_input_id = 14473 then
	sram_write <= x"22440220";
end if;
if first_state_sram_input_id = 14474 then
	sram_write <= x"C07C0068";
end if;
if first_state_sram_input_id = 14475 then
	sram_write <= x"D4264000";
end if;
if first_state_sram_input_id = 14476 then
	sram_write <= x"C03C0020";
end if;
if first_state_sram_input_id = 14477 then
	sram_write <= x"02220003";
end if;
if first_state_sram_input_id = 14478 then
	sram_write <= x"C05C0000";
end if;
if first_state_sram_input_id = 14479 then
	sram_write <= x"C4240000";
end if;
if first_state_sram_input_id = 14480 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 14481 then
	sram_write <= x"22220220";
end if;
if first_state_sram_input_id = 14482 then
	sram_write <= x"02220001";
end if;
if first_state_sram_input_id = 14483 then
	sram_write <= x"02600640";
end if;
if first_state_sram_input_id = 14484 then
	sram_write <= x"C0860000";
end if;
if first_state_sram_input_id = 14485 then
	sram_write <= x"C82000A8";
end if;
if first_state_sram_input_id = 14486 then
	sram_write <= x"C0A4001C";
end if;
if first_state_sram_input_id = 14487 then
	sram_write <= x"C84A0000";
end if;
if first_state_sram_input_id = 14488 then
	sram_write <= x"44224000";
end if;
if first_state_sram_input_id = 14489 then
	sram_write <= x"02A001D0";
end if;
if first_state_sram_input_id = 14490 then
	sram_write <= x"C0C40010";
end if;
if first_state_sram_input_id = 14491 then
	sram_write <= x"C84A0000";
end if;
if first_state_sram_input_id = 14492 then
	sram_write <= x"C86C0000";
end if;
if first_state_sram_input_id = 14493 then
	sram_write <= x"48446000";
end if;
if first_state_sram_input_id = 14494 then
	sram_write <= x"C86A0004";
end if;
if first_state_sram_input_id = 14495 then
	sram_write <= x"C88C0004";
end if;
if first_state_sram_input_id = 14496 then
	sram_write <= x"48668000";
end if;
if first_state_sram_input_id = 14497 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 14498 then
	sram_write <= x"C86A0008";
end if;
if first_state_sram_input_id = 14499 then
	sram_write <= x"C88C0008";
end if;
if first_state_sram_input_id = 14500 then
	sram_write <= x"48668000";
end if;
if first_state_sram_input_id = 14501 then
	sram_write <= x"40446000";
end if;
if first_state_sram_input_id = 14502 then
	sram_write <= x"C8600080";
end if;
if first_state_sram_input_id = 14503 then
	sram_write <= x"C0C40010";
end if;
if first_state_sram_input_id = 14504 then
	sram_write <= x"C88C0000";
end if;
if first_state_sram_input_id = 14505 then
	sram_write <= x"48868000";
end if;
if first_state_sram_input_id = 14506 then
	sram_write <= x"48884000";
end if;
if first_state_sram_input_id = 14507 then
	sram_write <= x"C8AA0000";
end if;
if first_state_sram_input_id = 14508 then
	sram_write <= x"4488A000";
end if;
if first_state_sram_input_id = 14509 then
	sram_write <= x"C0C40010";
end if;
if first_state_sram_input_id = 14510 then
	sram_write <= x"C8AC0004";
end if;
if first_state_sram_input_id = 14511 then
	sram_write <= x"48A6A000";
end if;
if first_state_sram_input_id = 14512 then
	sram_write <= x"48AA4000";
end if;
if first_state_sram_input_id = 14513 then
	sram_write <= x"C8CA0004";
end if;
if first_state_sram_input_id = 14514 then
	sram_write <= x"44AAC000";
end if;
if first_state_sram_input_id = 14515 then
	sram_write <= x"C0440010";
end if;
if first_state_sram_input_id = 14516 then
	sram_write <= x"C8C40008";
end if;
if first_state_sram_input_id = 14517 then
	sram_write <= x"4866C000";
end if;
if first_state_sram_input_id = 14518 then
	sram_write <= x"48464000";
end if;
if first_state_sram_input_id = 14519 then
	sram_write <= x"C86A0008";
end if;
if first_state_sram_input_id = 14520 then
	sram_write <= x"44446000";
end if;
if first_state_sram_input_id = 14521 then
	sram_write <= x"02400003";
end if;
if first_state_sram_input_id = 14522 then
	sram_write <= x"40600000";
end if;
if first_state_sram_input_id = 14523 then
	sram_write <= x"C47C0000";
end if;
if first_state_sram_input_id = 14524 then
	sram_write <= x"C49C0004";
end if;
if first_state_sram_input_id = 14525 then
	sram_write <= x"C43C0008";
end if;
if first_state_sram_input_id = 14526 then
	sram_write <= x"CC3C0010";
end if;
if first_state_sram_input_id = 14527 then
	sram_write <= x"CC5C0018";
end if;
if first_state_sram_input_id = 14528 then
	sram_write <= x"CCBC0020";
end if;
if first_state_sram_input_id = 14529 then
	sram_write <= x"CC9C0028";
end if;
if first_state_sram_input_id = 14530 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14531 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 14532 then
	sram_write <= x"40206000";
end if;
if first_state_sram_input_id = 14533 then
	sram_write <= x"03DC0038";
end if;
if first_state_sram_input_id = 14534 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14535 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14536 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 14537 then
	sram_write <= x"07DC0038";
end if;
if first_state_sram_input_id = 14538 then
	sram_write <= x"00420000";
end if;
if first_state_sram_input_id = 14539 then
	sram_write <= x"022000C4";
end if;
if first_state_sram_input_id = 14540 then
	sram_write <= x"C0620000";
end if;
if first_state_sram_input_id = 14541 then
	sram_write <= x"C43C0030";
end if;
if first_state_sram_input_id = 14542 then
	sram_write <= x"C45C0034";
end if;
if first_state_sram_input_id = 14543 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14544 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 14545 then
	sram_write <= x"03DC0040";
end if;
if first_state_sram_input_id = 14546 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14547 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14548 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 14549 then
	sram_write <= x"07DC0040";
end if;
if first_state_sram_input_id = 14550 then
	sram_write <= x"005A0000";
end if;
if first_state_sram_input_id = 14551 then
	sram_write <= x"03BA0008";
end if;
if first_state_sram_input_id = 14552 then
	sram_write <= x"C4240004";
end if;
if first_state_sram_input_id = 14553 then
	sram_write <= x"C07C0034";
end if;
if first_state_sram_input_id = 14554 then
	sram_write <= x"C4640000";
end if;
if first_state_sram_input_id = 14555 then
	sram_write <= x"C83C0028";
end if;
if first_state_sram_input_id = 14556 then
	sram_write <= x"CC260000";
end if;
if first_state_sram_input_id = 14557 then
	sram_write <= x"C83C0020";
end if;
if first_state_sram_input_id = 14558 then
	sram_write <= x"CC260004";
end if;
if first_state_sram_input_id = 14559 then
	sram_write <= x"C83C0018";
end if;
if first_state_sram_input_id = 14560 then
	sram_write <= x"CC260008";
end if;
if first_state_sram_input_id = 14561 then
	sram_write <= x"C09C0030";
end if;
if first_state_sram_input_id = 14562 then
	sram_write <= x"C0880000";
end if;
if first_state_sram_input_id = 14563 then
	sram_write <= x"06880001";
end if;
if first_state_sram_input_id = 14564 then
	sram_write <= x"C45C0038";
end if;
if first_state_sram_input_id = 14565 then
	sram_write <= x"8680E630";
end if;
if first_state_sram_input_id = 14566 then
	sram_write <= x"02A000C8";
end if;
if first_state_sram_input_id = 14567 then
	sram_write <= x"22C80220";
end if;
if first_state_sram_input_id = 14568 then
	sram_write <= x"D0CAC000";
end if;
if first_state_sram_input_id = 14569 then
	sram_write <= x"C0EC0004";
end if;
if first_state_sram_input_id = 14570 then
	sram_write <= x"03000001";
end if;
if first_state_sram_input_id = 14571 then
	sram_write <= x"C4BC003C";
end if;
if first_state_sram_input_id = 14572 then
	sram_write <= x"82F0E434";
end if;
if first_state_sram_input_id = 14573 then
	sram_write <= x"03000002";
end if;
if first_state_sram_input_id = 14574 then
	sram_write <= x"82F0E3F8";
end if;
if first_state_sram_input_id = 14575 then
	sram_write <= x"C43C0040";
end if;
if first_state_sram_input_id = 14576 then
	sram_write <= x"C49C0044";
end if;
if first_state_sram_input_id = 14577 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14578 then
	sram_write <= x"004C0000";
end if;
if first_state_sram_input_id = 14579 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 14580 then
	sram_write <= x"03DC0050";
end if;
if first_state_sram_input_id = 14581 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14582 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14583 then
	sram_write <= x"8200400C";
end if;
if first_state_sram_input_id = 14584 then
	sram_write <= x"07DC0050";
end if;
if first_state_sram_input_id = 14585 then
	sram_write <= x"C05C0044";
end if;
if first_state_sram_input_id = 14586 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 14587 then
	sram_write <= x"C09C0040";
end if;
if first_state_sram_input_id = 14588 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 14589 then
	sram_write <= x"8200E430";
end if;
if first_state_sram_input_id = 14590 then
	sram_write <= x"C43C0040";
end if;
if first_state_sram_input_id = 14591 then
	sram_write <= x"C49C0044";
end if;
if first_state_sram_input_id = 14592 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14593 then
	sram_write <= x"004C0000";
end if;
if first_state_sram_input_id = 14594 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 14595 then
	sram_write <= x"03DC0050";
end if;
if first_state_sram_input_id = 14596 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14597 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14598 then
	sram_write <= x"82003E98";
end if;
if first_state_sram_input_id = 14599 then
	sram_write <= x"07DC0050";
end if;
if first_state_sram_input_id = 14600 then
	sram_write <= x"C05C0044";
end if;
if first_state_sram_input_id = 14601 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 14602 then
	sram_write <= x"C09C0040";
end if;
if first_state_sram_input_id = 14603 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 14604 then
	sram_write <= x"8200E46C";
end if;
if first_state_sram_input_id = 14605 then
	sram_write <= x"C43C0040";
end if;
if first_state_sram_input_id = 14606 then
	sram_write <= x"C49C0044";
end if;
if first_state_sram_input_id = 14607 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14608 then
	sram_write <= x"004C0000";
end if;
if first_state_sram_input_id = 14609 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 14610 then
	sram_write <= x"03DC0050";
end if;
if first_state_sram_input_id = 14611 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14612 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14613 then
	sram_write <= x"82003CC4";
end if;
if first_state_sram_input_id = 14614 then
	sram_write <= x"07DC0050";
end if;
if first_state_sram_input_id = 14615 then
	sram_write <= x"C05C0044";
end if;
if first_state_sram_input_id = 14616 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 14617 then
	sram_write <= x"C09C0040";
end if;
if first_state_sram_input_id = 14618 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 14619 then
	sram_write <= x"06240001";
end if;
if first_state_sram_input_id = 14620 then
	sram_write <= x"8620E62C";
end if;
if first_state_sram_input_id = 14621 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 14622 then
	sram_write <= x"C07C003C";
end if;
if first_state_sram_input_id = 14623 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 14624 then
	sram_write <= x"C0A40004";
end if;
if first_state_sram_input_id = 14625 then
	sram_write <= x"02C00001";
end if;
if first_state_sram_input_id = 14626 then
	sram_write <= x"82ACE504";
end if;
if first_state_sram_input_id = 14627 then
	sram_write <= x"02C00002";
end if;
if first_state_sram_input_id = 14628 then
	sram_write <= x"82ACE4CC";
end if;
if first_state_sram_input_id = 14629 then
	sram_write <= x"C0BC0034";
end if;
if first_state_sram_input_id = 14630 then
	sram_write <= x"C43C0048";
end if;
if first_state_sram_input_id = 14631 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14632 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 14633 then
	sram_write <= x"03DC0054";
end if;
if first_state_sram_input_id = 14634 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14635 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14636 then
	sram_write <= x"8200400C";
end if;
if first_state_sram_input_id = 14637 then
	sram_write <= x"07DC0054";
end if;
if first_state_sram_input_id = 14638 then
	sram_write <= x"C05C0048";
end if;
if first_state_sram_input_id = 14639 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 14640 then
	sram_write <= x"C09C0040";
end if;
if first_state_sram_input_id = 14641 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 14642 then
	sram_write <= x"8200E500";
end if;
if first_state_sram_input_id = 14643 then
	sram_write <= x"C0BC0034";
end if;
if first_state_sram_input_id = 14644 then
	sram_write <= x"C43C0048";
end if;
if first_state_sram_input_id = 14645 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14646 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 14647 then
	sram_write <= x"03DC0054";
end if;
if first_state_sram_input_id = 14648 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14649 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14650 then
	sram_write <= x"82003E98";
end if;
if first_state_sram_input_id = 14651 then
	sram_write <= x"07DC0054";
end if;
if first_state_sram_input_id = 14652 then
	sram_write <= x"C05C0048";
end if;
if first_state_sram_input_id = 14653 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 14654 then
	sram_write <= x"C09C0040";
end if;
if first_state_sram_input_id = 14655 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 14656 then
	sram_write <= x"8200E538";
end if;
if first_state_sram_input_id = 14657 then
	sram_write <= x"C0BC0034";
end if;
if first_state_sram_input_id = 14658 then
	sram_write <= x"C43C0048";
end if;
if first_state_sram_input_id = 14659 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14660 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 14661 then
	sram_write <= x"03DC0054";
end if;
if first_state_sram_input_id = 14662 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14663 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14664 then
	sram_write <= x"82003CC4";
end if;
if first_state_sram_input_id = 14665 then
	sram_write <= x"07DC0054";
end if;
if first_state_sram_input_id = 14666 then
	sram_write <= x"C05C0048";
end if;
if first_state_sram_input_id = 14667 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 14668 then
	sram_write <= x"C09C0040";
end if;
if first_state_sram_input_id = 14669 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 14670 then
	sram_write <= x"06240001";
end if;
if first_state_sram_input_id = 14671 then
	sram_write <= x"8620E628";
end if;
if first_state_sram_input_id = 14672 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 14673 then
	sram_write <= x"C07C003C";
end if;
if first_state_sram_input_id = 14674 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 14675 then
	sram_write <= x"C0640004";
end if;
if first_state_sram_input_id = 14676 then
	sram_write <= x"02A00001";
end if;
if first_state_sram_input_id = 14677 then
	sram_write <= x"826AE5D0";
end if;
if first_state_sram_input_id = 14678 then
	sram_write <= x"02A00002";
end if;
if first_state_sram_input_id = 14679 then
	sram_write <= x"826AE598";
end if;
if first_state_sram_input_id = 14680 then
	sram_write <= x"C07C0034";
end if;
if first_state_sram_input_id = 14681 then
	sram_write <= x"C43C004C";
end if;
if first_state_sram_input_id = 14682 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14683 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 14684 then
	sram_write <= x"03DC0058";
end if;
if first_state_sram_input_id = 14685 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14686 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14687 then
	sram_write <= x"8200400C";
end if;
if first_state_sram_input_id = 14688 then
	sram_write <= x"07DC0058";
end if;
if first_state_sram_input_id = 14689 then
	sram_write <= x"C05C004C";
end if;
if first_state_sram_input_id = 14690 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 14691 then
	sram_write <= x"C09C0040";
end if;
if first_state_sram_input_id = 14692 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 14693 then
	sram_write <= x"8200E5CC";
end if;
if first_state_sram_input_id = 14694 then
	sram_write <= x"C07C0034";
end if;
if first_state_sram_input_id = 14695 then
	sram_write <= x"C43C004C";
end if;
if first_state_sram_input_id = 14696 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14697 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 14698 then
	sram_write <= x"03DC0058";
end if;
if first_state_sram_input_id = 14699 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14700 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14701 then
	sram_write <= x"82003E98";
end if;
if first_state_sram_input_id = 14702 then
	sram_write <= x"07DC0058";
end if;
if first_state_sram_input_id = 14703 then
	sram_write <= x"C05C004C";
end if;
if first_state_sram_input_id = 14704 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 14705 then
	sram_write <= x"C09C0040";
end if;
if first_state_sram_input_id = 14706 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 14707 then
	sram_write <= x"8200E604";
end if;
if first_state_sram_input_id = 14708 then
	sram_write <= x"C07C0034";
end if;
if first_state_sram_input_id = 14709 then
	sram_write <= x"C43C004C";
end if;
if first_state_sram_input_id = 14710 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14711 then
	sram_write <= x"00260000";
end if;
if first_state_sram_input_id = 14712 then
	sram_write <= x"03DC0058";
end if;
if first_state_sram_input_id = 14713 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14714 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14715 then
	sram_write <= x"82003CC4";
end if;
if first_state_sram_input_id = 14716 then
	sram_write <= x"07DC0058";
end if;
if first_state_sram_input_id = 14717 then
	sram_write <= x"C05C004C";
end if;
if first_state_sram_input_id = 14718 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 14719 then
	sram_write <= x"C09C0040";
end if;
if first_state_sram_input_id = 14720 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 14721 then
	sram_write <= x"06440001";
end if;
if first_state_sram_input_id = 14722 then
	sram_write <= x"C03C0038";
end if;
if first_state_sram_input_id = 14723 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14724 then
	sram_write <= x"03DC0058";
end if;
if first_state_sram_input_id = 14725 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14726 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14727 then
	sram_write <= x"820042A4";
end if;
if first_state_sram_input_id = 14728 then
	sram_write <= x"07DC0058";
end if;
if first_state_sram_input_id = 14729 then
	sram_write <= x"8200E628";
end if;
if first_state_sram_input_id = 14730 then
	sram_write <= x"8200E62C";
end if;
if first_state_sram_input_id = 14731 then
	sram_write <= x"8200E630";
end if;
if first_state_sram_input_id = 14732 then
	sram_write <= x"02200370";
end if;
if first_state_sram_input_id = 14733 then
	sram_write <= x"005A0000";
end if;
if first_state_sram_input_id = 14734 then
	sram_write <= x"03BA000C";
end if;
if first_state_sram_input_id = 14735 then
	sram_write <= x"C83C0010";
end if;
if first_state_sram_input_id = 14736 then
	sram_write <= x"CC240008";
end if;
if first_state_sram_input_id = 14737 then
	sram_write <= x"C07C0038";
end if;
if first_state_sram_input_id = 14738 then
	sram_write <= x"C4640004";
end if;
if first_state_sram_input_id = 14739 then
	sram_write <= x"C07C0008";
end if;
if first_state_sram_input_id = 14740 then
	sram_write <= x"C4640000";
end if;
if first_state_sram_input_id = 14741 then
	sram_write <= x"C07C0004";
end if;
if first_state_sram_input_id = 14742 then
	sram_write <= x"22860220";
end if;
if first_state_sram_input_id = 14743 then
	sram_write <= x"D4428000";
end if;
if first_state_sram_input_id = 14744 then
	sram_write <= x"02260001";
end if;
if first_state_sram_input_id = 14745 then
	sram_write <= x"C05C0000";
end if;
if first_state_sram_input_id = 14746 then
	sram_write <= x"C4240000";
end if;
if first_state_sram_input_id = 14747 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 14748 then
	sram_write <= x"026002F8";
end if;
if first_state_sram_input_id = 14749 then
	sram_write <= x"C4260000";
end if;
if first_state_sram_input_id = 14750 then
	sram_write <= x"C4460004";
end if;
if first_state_sram_input_id = 14751 then
	sram_write <= x"02800300";
end if;
if first_state_sram_input_id = 14752 then
	sram_write <= x"22A201A0";
end if;
if first_state_sram_input_id = 14753 then
	sram_write <= x"C4A80000";
end if;
if first_state_sram_input_id = 14754 then
	sram_write <= x"224401A0";
end if;
if first_state_sram_input_id = 14755 then
	sram_write <= x"C4480004";
end if;
if first_state_sram_input_id = 14756 then
	sram_write <= x"02400308";
end if;
if first_state_sram_input_id = 14757 then
	sram_write <= x"C8200004";
end if;
if first_state_sram_input_id = 14758 then
	sram_write <= x"58420000";
end if;
if first_state_sram_input_id = 14759 then
	sram_write <= x"C47C0000";
end if;
if first_state_sram_input_id = 14760 then
	sram_write <= x"C45C0004";
end if;
if first_state_sram_input_id = 14761 then
	sram_write <= x"CC3C0008";
end if;
if first_state_sram_input_id = 14762 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14763 then
	sram_write <= x"40204000";
end if;
if first_state_sram_input_id = 14764 then
	sram_write <= x"03DC0018";
end if;
if first_state_sram_input_id = 14765 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14766 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14767 then
	sram_write <= x"82000844";
end if;
if first_state_sram_input_id = 14768 then
	sram_write <= x"07DC0018";
end if;
if first_state_sram_input_id = 14769 then
	sram_write <= x"C85C0008";
end if;
if first_state_sram_input_id = 14770 then
	sram_write <= x"48242000";
end if;
if first_state_sram_input_id = 14771 then
	sram_write <= x"C03C0004";
end if;
if first_state_sram_input_id = 14772 then
	sram_write <= x"CC220000";
end if;
if first_state_sram_input_id = 14773 then
	sram_write <= x"C03C0000";
end if;
if first_state_sram_input_id = 14774 then
	sram_write <= x"C0420000";
end if;
if first_state_sram_input_id = 14775 then
	sram_write <= x"C45C0010";
end if;
if first_state_sram_input_id = 14776 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14777 then
	sram_write <= x"03DC001C";
end if;
if first_state_sram_input_id = 14778 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14779 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14780 then
	sram_write <= x"8200A47C";
end if;
if first_state_sram_input_id = 14781 then
	sram_write <= x"07DC001C";
end if;
if first_state_sram_input_id = 14782 then
	sram_write <= x"00420000";
end if;
if first_state_sram_input_id = 14783 then
	sram_write <= x"C03C0010";
end if;
if first_state_sram_input_id = 14784 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14785 then
	sram_write <= x"03DC001C";
end if;
if first_state_sram_input_id = 14786 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14787 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14788 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 14789 then
	sram_write <= x"07DC001C";
end if;
if first_state_sram_input_id = 14790 then
	sram_write <= x"C05C0000";
end if;
if first_state_sram_input_id = 14791 then
	sram_write <= x"C0640000";
end if;
if first_state_sram_input_id = 14792 then
	sram_write <= x"06660002";
end if;
if first_state_sram_input_id = 14793 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14794 then
	sram_write <= x"00460000";
end if;
if first_state_sram_input_id = 14795 then
	sram_write <= x"03DC001C";
end if;
if first_state_sram_input_id = 14796 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14797 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14798 then
	sram_write <= x"8200A914";
end if;
if first_state_sram_input_id = 14799 then
	sram_write <= x"07DC001C";
end if;
if first_state_sram_input_id = 14800 then
	sram_write <= x"C05C0000";
end if;
if first_state_sram_input_id = 14801 then
	sram_write <= x"C0640000";
end if;
if first_state_sram_input_id = 14802 then
	sram_write <= x"C43C0014";
end if;
if first_state_sram_input_id = 14803 then
	sram_write <= x"C47C0018";
end if;
if first_state_sram_input_id = 14804 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14805 then
	sram_write <= x"03DC0024";
end if;
if first_state_sram_input_id = 14806 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14807 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14808 then
	sram_write <= x"8200A47C";
end if;
if first_state_sram_input_id = 14809 then
	sram_write <= x"07DC0024";
end if;
if first_state_sram_input_id = 14810 then
	sram_write <= x"00420000";
end if;
if first_state_sram_input_id = 14811 then
	sram_write <= x"C03C0018";
end if;
if first_state_sram_input_id = 14812 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14813 then
	sram_write <= x"03DC0024";
end if;
if first_state_sram_input_id = 14814 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14815 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14816 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 14817 then
	sram_write <= x"07DC0024";
end if;
if first_state_sram_input_id = 14818 then
	sram_write <= x"C05C0000";
end if;
if first_state_sram_input_id = 14819 then
	sram_write <= x"C0640000";
end if;
if first_state_sram_input_id = 14820 then
	sram_write <= x"06660002";
end if;
if first_state_sram_input_id = 14821 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14822 then
	sram_write <= x"00460000";
end if;
if first_state_sram_input_id = 14823 then
	sram_write <= x"03DC0024";
end if;
if first_state_sram_input_id = 14824 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14825 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14826 then
	sram_write <= x"8200A914";
end if;
if first_state_sram_input_id = 14827 then
	sram_write <= x"07DC0024";
end if;
if first_state_sram_input_id = 14828 then
	sram_write <= x"C05C0000";
end if;
if first_state_sram_input_id = 14829 then
	sram_write <= x"C0640000";
end if;
if first_state_sram_input_id = 14830 then
	sram_write <= x"C43C001C";
end if;
if first_state_sram_input_id = 14831 then
	sram_write <= x"C47C0020";
end if;
if first_state_sram_input_id = 14832 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14833 then
	sram_write <= x"03DC002C";
end if;
if first_state_sram_input_id = 14834 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14835 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14836 then
	sram_write <= x"8200A47C";
end if;
if first_state_sram_input_id = 14837 then
	sram_write <= x"07DC002C";
end if;
if first_state_sram_input_id = 14838 then
	sram_write <= x"00420000";
end if;
if first_state_sram_input_id = 14839 then
	sram_write <= x"C03C0020";
end if;
if first_state_sram_input_id = 14840 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14841 then
	sram_write <= x"03DC002C";
end if;
if first_state_sram_input_id = 14842 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14843 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14844 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 14845 then
	sram_write <= x"07DC002C";
end if;
if first_state_sram_input_id = 14846 then
	sram_write <= x"C05C0000";
end if;
if first_state_sram_input_id = 14847 then
	sram_write <= x"C0640000";
end if;
if first_state_sram_input_id = 14848 then
	sram_write <= x"06660002";
end if;
if first_state_sram_input_id = 14849 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14850 then
	sram_write <= x"00460000";
end if;
if first_state_sram_input_id = 14851 then
	sram_write <= x"03DC002C";
end if;
if first_state_sram_input_id = 14852 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14853 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14854 then
	sram_write <= x"8200A914";
end if;
if first_state_sram_input_id = 14855 then
	sram_write <= x"07DC002C";
end if;
if first_state_sram_input_id = 14856 then
	sram_write <= x"C43C0024";
end if;
if first_state_sram_input_id = 14857 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14858 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 14859 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14860 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14861 then
	sram_write <= x"820016D4";
end if;
if first_state_sram_input_id = 14862 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 14863 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14864 then
	sram_write <= x"03DC0030";
end if;
if first_state_sram_input_id = 14865 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14866 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14867 then
	sram_write <= x"82001AB8";
end if;
if first_state_sram_input_id = 14868 then
	sram_write <= x"07DC0030";
end if;
if first_state_sram_input_id = 14869 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 14870 then
	sram_write <= x"C43C0028";
end if;
if first_state_sram_input_id = 14871 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14872 then
	sram_write <= x"03DC0034";
end if;
if first_state_sram_input_id = 14873 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14874 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14875 then
	sram_write <= x"82002384";
end if;
if first_state_sram_input_id = 14876 then
	sram_write <= x"07DC0034";
end if;
if first_state_sram_input_id = 14877 then
	sram_write <= x"8220E898";
end if;
if first_state_sram_input_id = 14878 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 14879 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14880 then
	sram_write <= x"03DC0034";
end if;
if first_state_sram_input_id = 14881 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14882 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14883 then
	sram_write <= x"82002930";
end if;
if first_state_sram_input_id = 14884 then
	sram_write <= x"07DC0034";
end if;
if first_state_sram_input_id = 14885 then
	sram_write <= x"8200E8A4";
end if;
if first_state_sram_input_id = 14886 then
	sram_write <= x"022000C4";
end if;
if first_state_sram_input_id = 14887 then
	sram_write <= x"C05C0028";
end if;
if first_state_sram_input_id = 14888 then
	sram_write <= x"C4420000";
end if;
if first_state_sram_input_id = 14889 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14890 then
	sram_write <= x"03DC0034";
end if;
if first_state_sram_input_id = 14891 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14892 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14893 then
	sram_write <= x"82000794";
end if;
if first_state_sram_input_id = 14894 then
	sram_write <= x"07DC0034";
end if;
if first_state_sram_input_id = 14895 then
	sram_write <= x"0240FFFF";
end if;
if first_state_sram_input_id = 14896 then
	sram_write <= x"8224E8F4";
end if;
if first_state_sram_input_id = 14897 then
	sram_write <= x"02400001";
end if;
if first_state_sram_input_id = 14898 then
	sram_write <= x"C43C002C";
end if;
if first_state_sram_input_id = 14899 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14900 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 14901 then
	sram_write <= x"03DC0038";
end if;
if first_state_sram_input_id = 14902 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14903 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14904 then
	sram_write <= x"82002A44";
end if;
if first_state_sram_input_id = 14905 then
	sram_write <= x"07DC0038";
end if;
if first_state_sram_input_id = 14906 then
	sram_write <= x"C05C002C";
end if;
if first_state_sram_input_id = 14907 then
	sram_write <= x"C4420000";
end if;
if first_state_sram_input_id = 14908 then
	sram_write <= x"8200E914";
end if;
if first_state_sram_input_id = 14909 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 14910 then
	sram_write <= x"0240FFFF";
end if;
if first_state_sram_input_id = 14911 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14912 then
	sram_write <= x"03DC0038";
end if;
if first_state_sram_input_id = 14913 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14914 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14915 then
	sram_write <= x"8200081C";
end if;
if first_state_sram_input_id = 14916 then
	sram_write <= x"07DC0038";
end if;
if first_state_sram_input_id = 14917 then
	sram_write <= x"C0420000";
end if;
if first_state_sram_input_id = 14918 then
	sram_write <= x"0260FFFF";
end if;
if first_state_sram_input_id = 14919 then
	sram_write <= x"8246E980";
end if;
if first_state_sram_input_id = 14920 then
	sram_write <= x"024001E0";
end if;
if first_state_sram_input_id = 14921 then
	sram_write <= x"C4240000";
end if;
if first_state_sram_input_id = 14922 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 14923 then
	sram_write <= x"C45C0030";
end if;
if first_state_sram_input_id = 14924 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14925 then
	sram_write <= x"03DC003C";
end if;
if first_state_sram_input_id = 14926 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14927 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14928 then
	sram_write <= x"82002A44";
end if;
if first_state_sram_input_id = 14929 then
	sram_write <= x"07DC003C";
end if;
if first_state_sram_input_id = 14930 then
	sram_write <= x"C0420000";
end if;
if first_state_sram_input_id = 14931 then
	sram_write <= x"0260FFFF";
end if;
if first_state_sram_input_id = 14932 then
	sram_write <= x"8246E97C";
end if;
if first_state_sram_input_id = 14933 then
	sram_write <= x"C05C0030";
end if;
if first_state_sram_input_id = 14934 then
	sram_write <= x"C4240004";
end if;
if first_state_sram_input_id = 14935 then
	sram_write <= x"02200002";
end if;
if first_state_sram_input_id = 14936 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14937 then
	sram_write <= x"03DC003C";
end if;
if first_state_sram_input_id = 14938 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14939 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14940 then
	sram_write <= x"82002E74";
end if;
if first_state_sram_input_id = 14941 then
	sram_write <= x"07DC003C";
end if;
if first_state_sram_input_id = 14942 then
	sram_write <= x"8200E97C";
end if;
if first_state_sram_input_id = 14943 then
	sram_write <= x"8200E980";
end if;
if first_state_sram_input_id = 14944 then
	sram_write <= x"022002A8";
end if;
if first_state_sram_input_id = 14945 then
	sram_write <= x"02400000";
end if;
if first_state_sram_input_id = 14946 then
	sram_write <= x"C43C0034";
end if;
if first_state_sram_input_id = 14947 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14948 then
	sram_write <= x"00240000";
end if;
if first_state_sram_input_id = 14949 then
	sram_write <= x"03DC0040";
end if;
if first_state_sram_input_id = 14950 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14951 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14952 then
	sram_write <= x"82002BEC";
end if;
if first_state_sram_input_id = 14953 then
	sram_write <= x"07DC0040";
end if;
if first_state_sram_input_id = 14954 then
	sram_write <= x"C05C0034";
end if;
if first_state_sram_input_id = 14955 then
	sram_write <= x"C4240000";
end if;
if first_state_sram_input_id = 14956 then
	sram_write <= x"02200050";
end if;
if first_state_sram_input_id = 14957 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14958 then
	sram_write <= x"03DC0040";
end if;
if first_state_sram_input_id = 14959 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14960 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14961 then
	sram_write <= x"8200078C";
end if;
if first_state_sram_input_id = 14962 then
	sram_write <= x"07DC0040";
end if;
if first_state_sram_input_id = 14963 then
	sram_write <= x"02200036";
end if;
if first_state_sram_input_id = 14964 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14965 then
	sram_write <= x"03DC0040";
end if;
if first_state_sram_input_id = 14966 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14967 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14968 then
	sram_write <= x"8200078C";
end if;
if first_state_sram_input_id = 14969 then
	sram_write <= x"07DC0040";
end if;
if first_state_sram_input_id = 14970 then
	sram_write <= x"0220000A";
end if;
if first_state_sram_input_id = 14971 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14972 then
	sram_write <= x"03DC0040";
end if;
if first_state_sram_input_id = 14973 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14974 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14975 then
	sram_write <= x"8200078C";
end if;
if first_state_sram_input_id = 14976 then
	sram_write <= x"07DC0040";
end if;
if first_state_sram_input_id = 14977 then
	sram_write <= x"02200031";
end if;
if first_state_sram_input_id = 14978 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14979 then
	sram_write <= x"03DC0040";
end if;
if first_state_sram_input_id = 14980 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14981 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14982 then
	sram_write <= x"8200078C";
end if;
if first_state_sram_input_id = 14983 then
	sram_write <= x"07DC0040";
end if;
if first_state_sram_input_id = 14984 then
	sram_write <= x"02200032";
end if;
if first_state_sram_input_id = 14985 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14986 then
	sram_write <= x"03DC0040";
end if;
if first_state_sram_input_id = 14987 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14988 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14989 then
	sram_write <= x"8200078C";
end if;
if first_state_sram_input_id = 14990 then
	sram_write <= x"07DC0040";
end if;
if first_state_sram_input_id = 14991 then
	sram_write <= x"02200038";
end if;
if first_state_sram_input_id = 14992 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 14993 then
	sram_write <= x"03DC0040";
end if;
if first_state_sram_input_id = 14994 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 14995 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 14996 then
	sram_write <= x"8200078C";
end if;
if first_state_sram_input_id = 14997 then
	sram_write <= x"07DC0040";
end if;
if first_state_sram_input_id = 14998 then
	sram_write <= x"02200020";
end if;
if first_state_sram_input_id = 14999 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 15000 then
	sram_write <= x"03DC0040";
end if;
if first_state_sram_input_id = 15001 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 15002 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 15003 then
	sram_write <= x"8200078C";
end if;
if first_state_sram_input_id = 15004 then
	sram_write <= x"07DC0040";
end if;
if first_state_sram_input_id = 15005 then
	sram_write <= x"02200031";
end if;
if first_state_sram_input_id = 15006 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 15007 then
	sram_write <= x"03DC0040";
end if;
if first_state_sram_input_id = 15008 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 15009 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 15010 then
	sram_write <= x"8200078C";
end if;
if first_state_sram_input_id = 15011 then
	sram_write <= x"07DC0040";
end if;
if first_state_sram_input_id = 15012 then
	sram_write <= x"02200032";
end if;
if first_state_sram_input_id = 15013 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 15014 then
	sram_write <= x"03DC0040";
end if;
if first_state_sram_input_id = 15015 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 15016 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 15017 then
	sram_write <= x"8200078C";
end if;
if first_state_sram_input_id = 15018 then
	sram_write <= x"07DC0040";
end if;
if first_state_sram_input_id = 15019 then
	sram_write <= x"02200038";
end if;
if first_state_sram_input_id = 15020 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 15021 then
	sram_write <= x"03DC0040";
end if;
if first_state_sram_input_id = 15022 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 15023 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 15024 then
	sram_write <= x"8200078C";
end if;
if first_state_sram_input_id = 15025 then
	sram_write <= x"07DC0040";
end if;
if first_state_sram_input_id = 15026 then
	sram_write <= x"0220000A";
end if;
if first_state_sram_input_id = 15027 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 15028 then
	sram_write <= x"03DC0040";
end if;
if first_state_sram_input_id = 15029 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 15030 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 15031 then
	sram_write <= x"8200078C";
end if;
if first_state_sram_input_id = 15032 then
	sram_write <= x"07DC0040";
end if;
if first_state_sram_input_id = 15033 then
	sram_write <= x"02200032";
end if;
if first_state_sram_input_id = 15034 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 15035 then
	sram_write <= x"03DC0040";
end if;
if first_state_sram_input_id = 15036 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 15037 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 15038 then
	sram_write <= x"8200078C";
end if;
if first_state_sram_input_id = 15039 then
	sram_write <= x"07DC0040";
end if;
if first_state_sram_input_id = 15040 then
	sram_write <= x"02200035";
end if;
if first_state_sram_input_id = 15041 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 15042 then
	sram_write <= x"03DC0040";
end if;
if first_state_sram_input_id = 15043 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 15044 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 15045 then
	sram_write <= x"8200078C";
end if;
if first_state_sram_input_id = 15046 then
	sram_write <= x"07DC0040";
end if;
if first_state_sram_input_id = 15047 then
	sram_write <= x"02200035";
end if;
if first_state_sram_input_id = 15048 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 15049 then
	sram_write <= x"03DC0040";
end if;
if first_state_sram_input_id = 15050 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 15051 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 15052 then
	sram_write <= x"8200078C";
end if;
if first_state_sram_input_id = 15053 then
	sram_write <= x"07DC0040";
end if;
if first_state_sram_input_id = 15054 then
	sram_write <= x"0220000A";
end if;
if first_state_sram_input_id = 15055 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 15056 then
	sram_write <= x"03DC0040";
end if;
if first_state_sram_input_id = 15057 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 15058 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 15059 then
	sram_write <= x"8200078C";
end if;
if first_state_sram_input_id = 15060 then
	sram_write <= x"07DC0040";
end if;
if first_state_sram_input_id = 15061 then
	sram_write <= x"02200004";
end if;
if first_state_sram_input_id = 15062 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 15063 then
	sram_write <= x"03DC0040";
end if;
if first_state_sram_input_id = 15064 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 15065 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 15066 then
	sram_write <= x"8200B92C";
end if;
if first_state_sram_input_id = 15067 then
	sram_write <= x"07DC0040";
end if;
if first_state_sram_input_id = 15068 then
	sram_write <= x"02200009";
end if;
if first_state_sram_input_id = 15069 then
	sram_write <= x"02400000";
end if;
if first_state_sram_input_id = 15070 then
	sram_write <= x"02600000";
end if;
if first_state_sram_input_id = 15071 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 15072 then
	sram_write <= x"03DC0040";
end if;
if first_state_sram_input_id = 15073 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 15074 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 15075 then
	sram_write <= x"8200B574";
end if;
if first_state_sram_input_id = 15076 then
	sram_write <= x"07DC0040";
end if;
if first_state_sram_input_id = 15077 then
	sram_write <= x"02200354";
end if;
if first_state_sram_input_id = 15078 then
	sram_write <= x"C0420010";
end if;
if first_state_sram_input_id = 15079 then
	sram_write <= x"C06401DC";
end if;
if first_state_sram_input_id = 15080 then
	sram_write <= x"028000C4";
end if;
if first_state_sram_input_id = 15081 then
	sram_write <= x"C0A80000";
end if;
if first_state_sram_input_id = 15082 then
	sram_write <= x"06AA0001";
end if;
if first_state_sram_input_id = 15083 then
	sram_write <= x"C49C0038";
end if;
if first_state_sram_input_id = 15084 then
	sram_write <= x"C43C003C";
end if;
if first_state_sram_input_id = 15085 then
	sram_write <= x"C45C0040";
end if;
if first_state_sram_input_id = 15086 then
	sram_write <= x"86A0EE78";
end if;
if first_state_sram_input_id = 15087 then
	sram_write <= x"02C000C8";
end if;
if first_state_sram_input_id = 15088 then
	sram_write <= x"22EA0220";
end if;
if first_state_sram_input_id = 15089 then
	sram_write <= x"D0ECE000";
end if;
if first_state_sram_input_id = 15090 then
	sram_write <= x"C1060004";
end if;
if first_state_sram_input_id = 15091 then
	sram_write <= x"C1260000";
end if;
if first_state_sram_input_id = 15092 then
	sram_write <= x"C14E0004";
end if;
if first_state_sram_input_id = 15093 then
	sram_write <= x"02800001";
end if;
if first_state_sram_input_id = 15094 then
	sram_write <= x"C47C0044";
end if;
if first_state_sram_input_id = 15095 then
	sram_write <= x"C4DC0048";
end if;
if first_state_sram_input_id = 15096 then
	sram_write <= x"8348EC64";
end if;
if first_state_sram_input_id = 15097 then
	sram_write <= x"02800002";
end if;
if first_state_sram_input_id = 15098 then
	sram_write <= x"8348EC28";
end if;
if first_state_sram_input_id = 15099 then
	sram_write <= x"C51C004C";
end if;
if first_state_sram_input_id = 15100 then
	sram_write <= x"C4BC0050";
end if;
if first_state_sram_input_id = 15101 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 15102 then
	sram_write <= x"004E0000";
end if;
if first_state_sram_input_id = 15103 then
	sram_write <= x"00320000";
end if;
if first_state_sram_input_id = 15104 then
	sram_write <= x"03DC005C";
end if;
if first_state_sram_input_id = 15105 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 15106 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 15107 then
	sram_write <= x"8200400C";
end if;
if first_state_sram_input_id = 15108 then
	sram_write <= x"07DC005C";
end if;
if first_state_sram_input_id = 15109 then
	sram_write <= x"C05C0050";
end if;
if first_state_sram_input_id = 15110 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 15111 then
	sram_write <= x"C09C004C";
end if;
if first_state_sram_input_id = 15112 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 15113 then
	sram_write <= x"8200EC60";
end if;
if first_state_sram_input_id = 15114 then
	sram_write <= x"C51C004C";
end if;
if first_state_sram_input_id = 15115 then
	sram_write <= x"C4BC0050";
end if;
if first_state_sram_input_id = 15116 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 15117 then
	sram_write <= x"004E0000";
end if;
if first_state_sram_input_id = 15118 then
	sram_write <= x"00320000";
end if;
if first_state_sram_input_id = 15119 then
	sram_write <= x"03DC005C";
end if;
if first_state_sram_input_id = 15120 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 15121 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 15122 then
	sram_write <= x"82003E98";
end if;
if first_state_sram_input_id = 15123 then
	sram_write <= x"07DC005C";
end if;
if first_state_sram_input_id = 15124 then
	sram_write <= x"C05C0050";
end if;
if first_state_sram_input_id = 15125 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 15126 then
	sram_write <= x"C09C004C";
end if;
if first_state_sram_input_id = 15127 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 15128 then
	sram_write <= x"8200EC9C";
end if;
if first_state_sram_input_id = 15129 then
	sram_write <= x"C51C004C";
end if;
if first_state_sram_input_id = 15130 then
	sram_write <= x"C4BC0050";
end if;
if first_state_sram_input_id = 15131 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 15132 then
	sram_write <= x"004E0000";
end if;
if first_state_sram_input_id = 15133 then
	sram_write <= x"00320000";
end if;
if first_state_sram_input_id = 15134 then
	sram_write <= x"03DC005C";
end if;
if first_state_sram_input_id = 15135 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 15136 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 15137 then
	sram_write <= x"82003CC4";
end if;
if first_state_sram_input_id = 15138 then
	sram_write <= x"07DC005C";
end if;
if first_state_sram_input_id = 15139 then
	sram_write <= x"C05C0050";
end if;
if first_state_sram_input_id = 15140 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 15141 then
	sram_write <= x"C09C004C";
end if;
if first_state_sram_input_id = 15142 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 15143 then
	sram_write <= x"06240001";
end if;
if first_state_sram_input_id = 15144 then
	sram_write <= x"8620EE74";
end if;
if first_state_sram_input_id = 15145 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 15146 then
	sram_write <= x"C07C0048";
end if;
if first_state_sram_input_id = 15147 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 15148 then
	sram_write <= x"C09C0044";
end if;
if first_state_sram_input_id = 15149 then
	sram_write <= x"C0A80004";
end if;
if first_state_sram_input_id = 15150 then
	sram_write <= x"C0C80000";
end if;
if first_state_sram_input_id = 15151 then
	sram_write <= x"C0E40004";
end if;
if first_state_sram_input_id = 15152 then
	sram_write <= x"03000001";
end if;
if first_state_sram_input_id = 15153 then
	sram_write <= x"82F0ED40";
end if;
if first_state_sram_input_id = 15154 then
	sram_write <= x"03000002";
end if;
if first_state_sram_input_id = 15155 then
	sram_write <= x"82F0ED08";
end if;
if first_state_sram_input_id = 15156 then
	sram_write <= x"C4BC0054";
end if;
if first_state_sram_input_id = 15157 then
	sram_write <= x"C43C0058";
end if;
if first_state_sram_input_id = 15158 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 15159 then
	sram_write <= x"002C0000";
end if;
if first_state_sram_input_id = 15160 then
	sram_write <= x"03DC0064";
end if;
if first_state_sram_input_id = 15161 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 15162 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 15163 then
	sram_write <= x"8200400C";
end if;
if first_state_sram_input_id = 15164 then
	sram_write <= x"07DC0064";
end if;
if first_state_sram_input_id = 15165 then
	sram_write <= x"C05C0058";
end if;
if first_state_sram_input_id = 15166 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 15167 then
	sram_write <= x"C09C0054";
end if;
if first_state_sram_input_id = 15168 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 15169 then
	sram_write <= x"8200ED3C";
end if;
if first_state_sram_input_id = 15170 then
	sram_write <= x"C4BC0054";
end if;
if first_state_sram_input_id = 15171 then
	sram_write <= x"C43C0058";
end if;
if first_state_sram_input_id = 15172 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 15173 then
	sram_write <= x"002C0000";
end if;
if first_state_sram_input_id = 15174 then
	sram_write <= x"03DC0064";
end if;
if first_state_sram_input_id = 15175 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 15176 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 15177 then
	sram_write <= x"82003E98";
end if;
if first_state_sram_input_id = 15178 then
	sram_write <= x"07DC0064";
end if;
if first_state_sram_input_id = 15179 then
	sram_write <= x"C05C0058";
end if;
if first_state_sram_input_id = 15180 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 15181 then
	sram_write <= x"C09C0054";
end if;
if first_state_sram_input_id = 15182 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 15183 then
	sram_write <= x"8200ED74";
end if;
if first_state_sram_input_id = 15184 then
	sram_write <= x"C4BC0054";
end if;
if first_state_sram_input_id = 15185 then
	sram_write <= x"C43C0058";
end if;
if first_state_sram_input_id = 15186 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 15187 then
	sram_write <= x"002C0000";
end if;
if first_state_sram_input_id = 15188 then
	sram_write <= x"03DC0064";
end if;
if first_state_sram_input_id = 15189 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 15190 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 15191 then
	sram_write <= x"82003CC4";
end if;
if first_state_sram_input_id = 15192 then
	sram_write <= x"07DC0064";
end if;
if first_state_sram_input_id = 15193 then
	sram_write <= x"C05C0058";
end if;
if first_state_sram_input_id = 15194 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 15195 then
	sram_write <= x"C09C0054";
end if;
if first_state_sram_input_id = 15196 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 15197 then
	sram_write <= x"06240001";
end if;
if first_state_sram_input_id = 15198 then
	sram_write <= x"8620EE70";
end if;
if first_state_sram_input_id = 15199 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 15200 then
	sram_write <= x"C07C0048";
end if;
if first_state_sram_input_id = 15201 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 15202 then
	sram_write <= x"C07C0044";
end if;
if first_state_sram_input_id = 15203 then
	sram_write <= x"C0860004";
end if;
if first_state_sram_input_id = 15204 then
	sram_write <= x"C0A60000";
end if;
if first_state_sram_input_id = 15205 then
	sram_write <= x"C0C40004";
end if;
if first_state_sram_input_id = 15206 then
	sram_write <= x"02E00001";
end if;
if first_state_sram_input_id = 15207 then
	sram_write <= x"82CEEE18";
end if;
if first_state_sram_input_id = 15208 then
	sram_write <= x"02E00002";
end if;
if first_state_sram_input_id = 15209 then
	sram_write <= x"82CEEDE0";
end if;
if first_state_sram_input_id = 15210 then
	sram_write <= x"C49C005C";
end if;
if first_state_sram_input_id = 15211 then
	sram_write <= x"C43C0060";
end if;
if first_state_sram_input_id = 15212 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 15213 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 15214 then
	sram_write <= x"03DC006C";
end if;
if first_state_sram_input_id = 15215 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 15216 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 15217 then
	sram_write <= x"8200400C";
end if;
if first_state_sram_input_id = 15218 then
	sram_write <= x"07DC006C";
end if;
if first_state_sram_input_id = 15219 then
	sram_write <= x"C05C0060";
end if;
if first_state_sram_input_id = 15220 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 15221 then
	sram_write <= x"C09C005C";
end if;
if first_state_sram_input_id = 15222 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 15223 then
	sram_write <= x"8200EE14";
end if;
if first_state_sram_input_id = 15224 then
	sram_write <= x"C49C005C";
end if;
if first_state_sram_input_id = 15225 then
	sram_write <= x"C43C0060";
end if;
if first_state_sram_input_id = 15226 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 15227 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 15228 then
	sram_write <= x"03DC006C";
end if;
if first_state_sram_input_id = 15229 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 15230 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 15231 then
	sram_write <= x"82003E98";
end if;
if first_state_sram_input_id = 15232 then
	sram_write <= x"07DC006C";
end if;
if first_state_sram_input_id = 15233 then
	sram_write <= x"C05C0060";
end if;
if first_state_sram_input_id = 15234 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 15235 then
	sram_write <= x"C09C005C";
end if;
if first_state_sram_input_id = 15236 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 15237 then
	sram_write <= x"8200EE4C";
end if;
if first_state_sram_input_id = 15238 then
	sram_write <= x"C49C005C";
end if;
if first_state_sram_input_id = 15239 then
	sram_write <= x"C43C0060";
end if;
if first_state_sram_input_id = 15240 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 15241 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 15242 then
	sram_write <= x"03DC006C";
end if;
if first_state_sram_input_id = 15243 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 15244 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 15245 then
	sram_write <= x"82003CC4";
end if;
if first_state_sram_input_id = 15246 then
	sram_write <= x"07DC006C";
end if;
if first_state_sram_input_id = 15247 then
	sram_write <= x"C05C0060";
end if;
if first_state_sram_input_id = 15248 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 15249 then
	sram_write <= x"C09C005C";
end if;
if first_state_sram_input_id = 15250 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 15251 then
	sram_write <= x"06440001";
end if;
if first_state_sram_input_id = 15252 then
	sram_write <= x"C03C0044";
end if;
if first_state_sram_input_id = 15253 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 15254 then
	sram_write <= x"03DC006C";
end if;
if first_state_sram_input_id = 15255 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 15256 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 15257 then
	sram_write <= x"820042A4";
end if;
if first_state_sram_input_id = 15258 then
	sram_write <= x"07DC006C";
end if;
if first_state_sram_input_id = 15259 then
	sram_write <= x"8200EE70";
end if;
if first_state_sram_input_id = 15260 then
	sram_write <= x"8200EE74";
end if;
if first_state_sram_input_id = 15261 then
	sram_write <= x"8200EE78";
end if;
if first_state_sram_input_id = 15262 then
	sram_write <= x"02400076";
end if;
if first_state_sram_input_id = 15263 then
	sram_write <= x"C03C0040";
end if;
if first_state_sram_input_id = 15264 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 15265 then
	sram_write <= x"03DC006C";
end if;
if first_state_sram_input_id = 15266 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 15267 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 15268 then
	sram_write <= x"8200BD10";
end if;
if first_state_sram_input_id = 15269 then
	sram_write <= x"07DC006C";
end if;
if first_state_sram_input_id = 15270 then
	sram_write <= x"C03C003C";
end if;
if first_state_sram_input_id = 15271 then
	sram_write <= x"C022000C";
end if;
if first_state_sram_input_id = 15272 then
	sram_write <= x"02400077";
end if;
if first_state_sram_input_id = 15273 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 15274 then
	sram_write <= x"03DC006C";
end if;
if first_state_sram_input_id = 15275 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 15276 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 15277 then
	sram_write <= x"8200BD10";
end if;
if first_state_sram_input_id = 15278 then
	sram_write <= x"07DC006C";
end if;
if first_state_sram_input_id = 15279 then
	sram_write <= x"02200002";
end if;
if first_state_sram_input_id = 15280 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 15281 then
	sram_write <= x"03DC006C";
end if;
if first_state_sram_input_id = 15282 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 15283 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 15284 then
	sram_write <= x"8200C714";
end if;
if first_state_sram_input_id = 15285 then
	sram_write <= x"07DC006C";
end if;
if first_state_sram_input_id = 15286 then
	sram_write <= x"02200368";
end if;
if first_state_sram_input_id = 15287 then
	sram_write <= x"C0420000";
end if;
if first_state_sram_input_id = 15288 then
	sram_write <= x"026001D0";
end if;
if first_state_sram_input_id = 15289 then
	sram_write <= x"C8260000";
end if;
if first_state_sram_input_id = 15290 then
	sram_write <= x"CC240000";
end if;
if first_state_sram_input_id = 15291 then
	sram_write <= x"C8260004";
end if;
if first_state_sram_input_id = 15292 then
	sram_write <= x"CC240004";
end if;
if first_state_sram_input_id = 15293 then
	sram_write <= x"C8260008";
end if;
if first_state_sram_input_id = 15294 then
	sram_write <= x"CC240008";
end if;
if first_state_sram_input_id = 15295 then
	sram_write <= x"C05C0038";
end if;
if first_state_sram_input_id = 15296 then
	sram_write <= x"C0640000";
end if;
if first_state_sram_input_id = 15297 then
	sram_write <= x"06660001";
end if;
if first_state_sram_input_id = 15298 then
	sram_write <= x"8660F0EC";
end if;
if first_state_sram_input_id = 15299 then
	sram_write <= x"028000C8";
end if;
if first_state_sram_input_id = 15300 then
	sram_write <= x"22A60220";
end if;
if first_state_sram_input_id = 15301 then
	sram_write <= x"D0A8A000";
end if;
if first_state_sram_input_id = 15302 then
	sram_write <= x"C0C20004";
end if;
if first_state_sram_input_id = 15303 then
	sram_write <= x"C0E20000";
end if;
if first_state_sram_input_id = 15304 then
	sram_write <= x"C10A0004";
end if;
if first_state_sram_input_id = 15305 then
	sram_write <= x"03200001";
end if;
if first_state_sram_input_id = 15306 then
	sram_write <= x"C43C0064";
end if;
if first_state_sram_input_id = 15307 then
	sram_write <= x"C49C0068";
end if;
if first_state_sram_input_id = 15308 then
	sram_write <= x"8312EFB4";
end if;
if first_state_sram_input_id = 15309 then
	sram_write <= x"03200002";
end if;
if first_state_sram_input_id = 15310 then
	sram_write <= x"8312EF78";
end if;
if first_state_sram_input_id = 15311 then
	sram_write <= x"C4DC006C";
end if;
if first_state_sram_input_id = 15312 then
	sram_write <= x"C47C0070";
end if;
if first_state_sram_input_id = 15313 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 15314 then
	sram_write <= x"004A0000";
end if;
if first_state_sram_input_id = 15315 then
	sram_write <= x"002E0000";
end if;
if first_state_sram_input_id = 15316 then
	sram_write <= x"03DC007C";
end if;
if first_state_sram_input_id = 15317 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 15318 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 15319 then
	sram_write <= x"8200400C";
end if;
if first_state_sram_input_id = 15320 then
	sram_write <= x"07DC007C";
end if;
if first_state_sram_input_id = 15321 then
	sram_write <= x"C05C0070";
end if;
if first_state_sram_input_id = 15322 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 15323 then
	sram_write <= x"C09C006C";
end if;
if first_state_sram_input_id = 15324 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 15325 then
	sram_write <= x"8200EFB0";
end if;
if first_state_sram_input_id = 15326 then
	sram_write <= x"C4DC006C";
end if;
if first_state_sram_input_id = 15327 then
	sram_write <= x"C47C0070";
end if;
if first_state_sram_input_id = 15328 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 15329 then
	sram_write <= x"004A0000";
end if;
if first_state_sram_input_id = 15330 then
	sram_write <= x"002E0000";
end if;
if first_state_sram_input_id = 15331 then
	sram_write <= x"03DC007C";
end if;
if first_state_sram_input_id = 15332 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 15333 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 15334 then
	sram_write <= x"82003E98";
end if;
if first_state_sram_input_id = 15335 then
	sram_write <= x"07DC007C";
end if;
if first_state_sram_input_id = 15336 then
	sram_write <= x"C05C0070";
end if;
if first_state_sram_input_id = 15337 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 15338 then
	sram_write <= x"C09C006C";
end if;
if first_state_sram_input_id = 15339 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 15340 then
	sram_write <= x"8200EFEC";
end if;
if first_state_sram_input_id = 15341 then
	sram_write <= x"C4DC006C";
end if;
if first_state_sram_input_id = 15342 then
	sram_write <= x"C47C0070";
end if;
if first_state_sram_input_id = 15343 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 15344 then
	sram_write <= x"004A0000";
end if;
if first_state_sram_input_id = 15345 then
	sram_write <= x"002E0000";
end if;
if first_state_sram_input_id = 15346 then
	sram_write <= x"03DC007C";
end if;
if first_state_sram_input_id = 15347 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 15348 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 15349 then
	sram_write <= x"82003CC4";
end if;
if first_state_sram_input_id = 15350 then
	sram_write <= x"07DC007C";
end if;
if first_state_sram_input_id = 15351 then
	sram_write <= x"C05C0070";
end if;
if first_state_sram_input_id = 15352 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 15353 then
	sram_write <= x"C09C006C";
end if;
if first_state_sram_input_id = 15354 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 15355 then
	sram_write <= x"06240001";
end if;
if first_state_sram_input_id = 15356 then
	sram_write <= x"8620F0E8";
end if;
if first_state_sram_input_id = 15357 then
	sram_write <= x"22420220";
end if;
if first_state_sram_input_id = 15358 then
	sram_write <= x"C07C0068";
end if;
if first_state_sram_input_id = 15359 then
	sram_write <= x"D0464000";
end if;
if first_state_sram_input_id = 15360 then
	sram_write <= x"C07C0064";
end if;
if first_state_sram_input_id = 15361 then
	sram_write <= x"C0860004";
end if;
if first_state_sram_input_id = 15362 then
	sram_write <= x"C0A60000";
end if;
if first_state_sram_input_id = 15363 then
	sram_write <= x"C0C40004";
end if;
if first_state_sram_input_id = 15364 then
	sram_write <= x"02E00001";
end if;
if first_state_sram_input_id = 15365 then
	sram_write <= x"82CEF090";
end if;
if first_state_sram_input_id = 15366 then
	sram_write <= x"02E00002";
end if;
if first_state_sram_input_id = 15367 then
	sram_write <= x"82CEF058";
end if;
if first_state_sram_input_id = 15368 then
	sram_write <= x"C49C0074";
end if;
if first_state_sram_input_id = 15369 then
	sram_write <= x"C43C0078";
end if;
if first_state_sram_input_id = 15370 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 15371 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 15372 then
	sram_write <= x"03DC0084";
end if;
if first_state_sram_input_id = 15373 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 15374 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 15375 then
	sram_write <= x"8200400C";
end if;
if first_state_sram_input_id = 15376 then
	sram_write <= x"07DC0084";
end if;
if first_state_sram_input_id = 15377 then
	sram_write <= x"C05C0078";
end if;
if first_state_sram_input_id = 15378 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 15379 then
	sram_write <= x"C09C0074";
end if;
if first_state_sram_input_id = 15380 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 15381 then
	sram_write <= x"8200F08C";
end if;
if first_state_sram_input_id = 15382 then
	sram_write <= x"C49C0074";
end if;
if first_state_sram_input_id = 15383 then
	sram_write <= x"C43C0078";
end if;
if first_state_sram_input_id = 15384 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 15385 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 15386 then
	sram_write <= x"03DC0084";
end if;
if first_state_sram_input_id = 15387 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 15388 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 15389 then
	sram_write <= x"82003E98";
end if;
if first_state_sram_input_id = 15390 then
	sram_write <= x"07DC0084";
end if;
if first_state_sram_input_id = 15391 then
	sram_write <= x"C05C0078";
end if;
if first_state_sram_input_id = 15392 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 15393 then
	sram_write <= x"C09C0074";
end if;
if first_state_sram_input_id = 15394 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 15395 then
	sram_write <= x"8200F0C4";
end if;
if first_state_sram_input_id = 15396 then
	sram_write <= x"C49C0074";
end if;
if first_state_sram_input_id = 15397 then
	sram_write <= x"C43C0078";
end if;
if first_state_sram_input_id = 15398 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 15399 then
	sram_write <= x"002A0000";
end if;
if first_state_sram_input_id = 15400 then
	sram_write <= x"03DC0084";
end if;
if first_state_sram_input_id = 15401 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 15402 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 15403 then
	sram_write <= x"82003CC4";
end if;
if first_state_sram_input_id = 15404 then
	sram_write <= x"07DC0084";
end if;
if first_state_sram_input_id = 15405 then
	sram_write <= x"C05C0078";
end if;
if first_state_sram_input_id = 15406 then
	sram_write <= x"22640220";
end if;
if first_state_sram_input_id = 15407 then
	sram_write <= x"C09C0074";
end if;
if first_state_sram_input_id = 15408 then
	sram_write <= x"D4286000";
end if;
if first_state_sram_input_id = 15409 then
	sram_write <= x"06440001";
end if;
if first_state_sram_input_id = 15410 then
	sram_write <= x"C03C0064";
end if;
if first_state_sram_input_id = 15411 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 15412 then
	sram_write <= x"03DC0084";
end if;
if first_state_sram_input_id = 15413 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 15414 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 15415 then
	sram_write <= x"820042A4";
end if;
if first_state_sram_input_id = 15416 then
	sram_write <= x"07DC0084";
end if;
if first_state_sram_input_id = 15417 then
	sram_write <= x"8200F0E8";
end if;
if first_state_sram_input_id = 15418 then
	sram_write <= x"8200F0EC";
end if;
if first_state_sram_input_id = 15419 then
	sram_write <= x"C03C0038";
end if;
if first_state_sram_input_id = 15420 then
	sram_write <= x"C0220000";
end if;
if first_state_sram_input_id = 15421 then
	sram_write <= x"06220001";
end if;
if first_state_sram_input_id = 15422 then
	sram_write <= x"8620F17C";
end if;
if first_state_sram_input_id = 15423 then
	sram_write <= x"024000C8";
end if;
if first_state_sram_input_id = 15424 then
	sram_write <= x"22620220";
end if;
if first_state_sram_input_id = 15425 then
	sram_write <= x"D0446000";
end if;
if first_state_sram_input_id = 15426 then
	sram_write <= x"C0640008";
end if;
if first_state_sram_input_id = 15427 then
	sram_write <= x"02800002";
end if;
if first_state_sram_input_id = 15428 then
	sram_write <= x"8268F118";
end if;
if first_state_sram_input_id = 15429 then
	sram_write <= x"8200F178";
end if;
if first_state_sram_input_id = 15430 then
	sram_write <= x"C064001C";
end if;
if first_state_sram_input_id = 15431 then
	sram_write <= x"C8260000";
end if;
if first_state_sram_input_id = 15432 then
	sram_write <= x"C84000A8";
end if;
if first_state_sram_input_id = 15433 then
	sram_write <= x"8E24F12C";
end if;
if first_state_sram_input_id = 15434 then
	sram_write <= x"8200F178";
end if;
if first_state_sram_input_id = 15435 then
	sram_write <= x"C0640004";
end if;
if first_state_sram_input_id = 15436 then
	sram_write <= x"02800001";
end if;
if first_state_sram_input_id = 15437 then
	sram_write <= x"8268F160";
end if;
if first_state_sram_input_id = 15438 then
	sram_write <= x"02800002";
end if;
if first_state_sram_input_id = 15439 then
	sram_write <= x"8268F144";
end if;
if first_state_sram_input_id = 15440 then
	sram_write <= x"8200F15C";
end if;
if first_state_sram_input_id = 15441 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 15442 then
	sram_write <= x"03DC0084";
end if;
if first_state_sram_input_id = 15443 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 15444 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 15445 then
	sram_write <= x"8200E244";
end if;
if first_state_sram_input_id = 15446 then
	sram_write <= x"07DC0084";
end if;
if first_state_sram_input_id = 15447 then
	sram_write <= x"8200F178";
end if;
if first_state_sram_input_id = 15448 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 15449 then
	sram_write <= x"03DC0084";
end if;
if first_state_sram_input_id = 15450 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 15451 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 15452 then
	sram_write <= x"8200D764";
end if;
if first_state_sram_input_id = 15453 then
	sram_write <= x"07DC0084";
end if;
if first_state_sram_input_id = 15454 then
	sram_write <= x"8200F17C";
end if;
if first_state_sram_input_id = 15455 then
	sram_write <= x"02400000";
end if;
if first_state_sram_input_id = 15456 then
	sram_write <= x"02600000";
end if;
if first_state_sram_input_id = 15457 then
	sram_write <= x"C03C001C";
end if;
if first_state_sram_input_id = 15458 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 15459 then
	sram_write <= x"03DC0084";
end if;
if first_state_sram_input_id = 15460 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 15461 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 15462 then
	sram_write <= x"82009C08";
end if;
if first_state_sram_input_id = 15463 then
	sram_write <= x"07DC0084";
end if;
if first_state_sram_input_id = 15464 then
	sram_write <= x"02400000";
end if;
if first_state_sram_input_id = 15465 then
	sram_write <= x"02600002";
end if;
if first_state_sram_input_id = 15466 then
	sram_write <= x"C03C0000";
end if;
if first_state_sram_input_id = 15467 then
	sram_write <= x"C0820004";
end if;
if first_state_sram_input_id = 15468 then
	sram_write <= x"8608F1B8";
end if;
if first_state_sram_input_id = 15469 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 15470 then
	sram_write <= x"C0220004";
end if;
if first_state_sram_input_id = 15471 then
	sram_write <= x"06220001";
end if;
if first_state_sram_input_id = 15472 then
	sram_write <= x"C45C007C";
end if;
if first_state_sram_input_id = 15473 then
	sram_write <= x"8602F1CC";
end if;
if first_state_sram_input_id = 15474 then
	sram_write <= x"8200F1F4";
end if;
if first_state_sram_input_id = 15475 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 15476 then
	sram_write <= x"C09C0024";
end if;
if first_state_sram_input_id = 15477 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 15478 then
	sram_write <= x"00420000";
end if;
if first_state_sram_input_id = 15479 then
	sram_write <= x"00280000";
end if;
if first_state_sram_input_id = 15480 then
	sram_write <= x"03DC0088";
end if;
if first_state_sram_input_id = 15481 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 15482 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 15483 then
	sram_write <= x"82009C08";
end if;
if first_state_sram_input_id = 15484 then
	sram_write <= x"07DC0088";
end if;
if first_state_sram_input_id = 15485 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 15486 then
	sram_write <= x"C05C007C";
end if;
if first_state_sram_input_id = 15487 then
	sram_write <= x"C07C0014";
end if;
if first_state_sram_input_id = 15488 then
	sram_write <= x"C09C001C";
end if;
if first_state_sram_input_id = 15489 then
	sram_write <= x"C0BC0024";
end if;
if first_state_sram_input_id = 15490 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 15491 then
	sram_write <= x"03DC0088";
end if;
if first_state_sram_input_id = 15492 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 15493 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 15494 then
	sram_write <= x"82009C7C";
end if;
if first_state_sram_input_id = 15495 then
	sram_write <= x"07DC0088";
end if;
if first_state_sram_input_id = 15496 then
	sram_write <= x"02200001";
end if;
if first_state_sram_input_id = 15497 then
	sram_write <= x"02A00004";
end if;
if first_state_sram_input_id = 15498 then
	sram_write <= x"C05C001C";
end if;
if first_state_sram_input_id = 15499 then
	sram_write <= x"C07C0024";
end if;
if first_state_sram_input_id = 15500 then
	sram_write <= x"C09C0014";
end if;
if first_state_sram_input_id = 15501 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 15502 then
	sram_write <= x"03DC0088";
end if;
if first_state_sram_input_id = 15503 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 15504 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 15505 then
	sram_write <= x"8200A164";
end if;
if first_state_sram_input_id = 15506 then
	sram_write <= x"07DC0088";
end if;
if first_state_sram_input_id = 15507 then
	sram_write <= x"C1FDFFFC";
end if;
if first_state_sram_input_id = 15508 then
	sram_write <= x"03DC0004";
end if;
if first_state_sram_input_id = 15509 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 15510 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 15511 then
	sram_write <= x"82000644";
end if;
if first_state_sram_input_id = 15512 then
	sram_write <= x"07DC0004";
end if;
if first_state_sram_input_id = 15513 then
	sram_write <= x"02200080";
end if;
if first_state_sram_input_id = 15514 then
	sram_write <= x"02400080";
end if;
if first_state_sram_input_id = 15515 then
	sram_write <= x"C17DFFFC";
end if;
if first_state_sram_input_id = 15516 then
	sram_write <= x"03DC0008";
end if;
if first_state_sram_input_id = 15517 then
	sram_write <= x"037E000C";
end if;
if first_state_sram_input_id = 15518 then
	sram_write <= x"C57DFFFC";
end if;
if first_state_sram_input_id = 15519 then
	sram_write <= x"8200E670";
end if;
if first_state_sram_input_id = 15520 then
	sram_write <= x"07DC0008";
end if;
if first_state_sram_input_id = 15521 then
	sram_write <= x"02200000";
end if;
if first_state_sram_input_id = 15522 then
	sram_write <= x"8001E000";
end if;
            else
              sram_go <= '0';
            end if;
          else
            sram_go <= '0';
            top_state <= "001";
          end if;
        else
          if (first_state_write_wait = 5) then
            if first_state_sram_input_id = 15522 then
              first_state_sram_input_id <= x"55555";
            else
              first_state_sram_input_id <= first_state_sram_input_id + 1;
            end if;
          end if;
          if (first_state_write_wait > 0) then
            first_state_write_wait <= first_state_write_wait - 1;
          end if;
          sram_go <= '0';
        end if;
      end if;
      if top_state = "001" then
        --Input Wait
        if exok_from_read = '1' then
          exok <= '1';
          top_state <= "010";
          --if u232c_busy = '0' then
          --  u232c_data_reg <= x"000000" & debug_otpt_inputc;
          --  u232c_showtype <= "000";
          --  u232c_go <= '1';
          --else
          --  u232c_go <= '0';
          --end if;
        end if;
        if sram_busy = '0' then
          if inputc_write_ok = '1' then
            sram_go <= '1';
            --write
            sram_inst_type <= '1';
            sram_addr <= inputc_write_addr;
            sram_write <= inputc_write_value;
            debug_saved_value <= inputc_write_value;
            sigcount <= x"8";
            if u232c_busy = '0' then
              u232c_data_reg <= inputc_write_value;
              u232c_showtype <= "000";
              u232c_go <= '1';
            else
              u232c_go <= '0';
            end if;
          else
            u232c_go <= '0';
            sram_go <= '0';
          end if;
        else
          u232c_go <= '0';
          sram_go <= '0';
        end if;
      end if;
      if top_state = "010" then
        --Execution
        if u232c_busy = '0' then
          u232c_data_reg <= debug_otpt;
          u232c_showtype <= debug_otpt_code;
          u232c_go <= debug_otpt_signal;
        else
          u232c_go <= '0';
        end if;
        -- 垂れ流し
        core_sram_read <= sram_read;
        if sram_busy = '0' then
          if core_sram_go = '1' then
            sram_go <= '1';
            if core_sram_inst_type = '0' then
              --read
              sram_inst_type <= '0';
              sram_addr <= core_sram_addr;
            else
              --write
              sram_inst_type <= '1';
              sram_addr <= core_sram_addr;
              sram_write <= core_sram_write;
            end if;
          else
            sram_go <= '0';
          end if;
        else
          sram_go <= '0';
        end if;
      end if;
    end if;
  end process;
end cpu_top;

