-- CORE
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity core is
  Port (
    clk : in std_logic;
    execute_ok : in std_logic;
    ostate : out std_logic_vector(7 downto 0);
    sram_go : out std_logic := '0';
    sram_inst_type : out std_logic;
    sram_addr : out std_logic_vector(19 downto 0);
    sram_read : in std_logic_vector(31 downto 0);
    sram_write : out std_logic_vector(31 downto 0);
    debug_otpt : out std_logic_vector(7 downto 0);
    debug_otpt_signal : out std_logic := '0';
    waitwrite_from_parent : in std_logic_vector(19 downto 0);
    read_signal : out std_logic := '0'
  );
end core;

architecture cocore of core is
--components
  component alu Port (
    clk : in std_logic;
    opc_alu : in std_logic_vector(6 downto 0);
    reg_in_a : in std_logic_vector(31 downto 0);
    reg_in_b : in std_logic_vector(31 downto 0);
    reg_out : out std_logic_vector(31 downto 0);
    shift_dir : in std_logic;
    shift_type : in std_logic_vector(1 downto 0);
    shift_go : in std_logic
  );
  end component;
  component compr Port (
    clk : in std_logic;
    opc_compr : in std_logic_vector(6 downto 0);
    reg_in_a : in std_logic_vector(31 downto 0);
    reg_in_b : in std_logic_vector(31 downto 0);
    cond_out : out std_logic
  );
  end component;
  component fpu_man Port (
    clk : in std_logic;
    opc_fpu : in std_logic_vector(6 downto 0);
    reg_in_a : in std_logic_vector(31 downto 0);
    reg_in_b : in std_logic_vector(31 downto 0);
    reg_out : out std_logic_vector(31 downto 0)
  );
  end component;
  -- registers
  type registers is array (15 downto 0) of std_logic_vector (31 downto 0);
  -- rg (13) : hp ,rg (14) : sp ,rg (15) : pc ,
  signal rg : registers := (13 => x"00155554",14 => x"002AAAA8",others => (others => '0'));
  signal fp : registers := (others => (others => '0'));

-- signals
  signal state : std_logic_vector(7 downto 0) := x"00";
  signal phase : std_logic_vector(2 downto 0) := "111";
    --phase: active phase (without pipelines)
  signal cond_new_pc : std_logic_vector(31 downto 0) := x"00000000";
  signal opccode_alu : std_logic_vector(6 downto 0);
  signal reg_in_a : std_logic_vector(31 downto 0);
  signal reg_in_b : std_logic_vector(31 downto 0);
  signal reg_out : std_logic_vector(31 downto 0);
  signal shift_dir : std_logic;
  signal shift_type : std_logic_vector(1 downto 0);
  signal shift_go : std_logic := '0';
  signal opccode_fpu : std_logic_vector(6 downto 0);
  signal reg_in_a_fpu : std_logic_vector(31 downto 0);
  signal reg_in_b_fpu : std_logic_vector(31 downto 0);
  signal reg_out_fpu : std_logic_vector(31 downto 0);
  signal opccode_compr : std_logic_vector(6 downto 0);
  signal reg_in_a_compr : std_logic_vector(31 downto 0);
  signal reg_in_b_compr : std_logic_vector(31 downto 0);
  signal cond_out_compr : std_logic;
  signal dest_reg : std_logic_vector(3 downto 0);
  signal loaded_srca : std_logic_vector(31 downto 0);
  signal loaded_srcb : std_logic_vector(31 downto 0);
  signal loaded_newpc : std_logic_vector(31 downto 0);
  signal read_index : std_logic_vector(19 downto 0) := x"00000";
  signal waitwriting : std_logic := '0';
  type cache_array is array(16383 downto 0) of std_logic_vector(31 downto 0);
  signal cache_inst : cache_array := (x"8200F250",x"43000000",x"BDCCCCCD",x"3F666666",x"3E4CCCCD",x"C3160000",x"43160000",x"3DCCCCCD",x"C0000000",x"43800000",x"4CBEBC20",x"4E6E6B28",x"41A00000",x"3D4CCCCD",x"3E800000",x"41200000",x"3E99999A",x"437F0000",x"3E19999A",x"41700000",x"40490FDC",x"41F00000",x"3C75989E",x"3F6DA101",x"3C8F53C5",x"3E0E9468",x"3CF30835",x"38D1B717",x"BDCCCCCD",x"3C23D70A",x"BE4CCCCD",x"BF800000",x"40000000",x"C3480000",x"43480000",x"3C8EF998",x"C0C90FDA",x"00000000",x"40C90FDA",x"3AB39192",x"3D2AA7DF",x"3F000000",x"3F800000",x"394D8559",x"3C088723",x"3E2AAAC1",x"3F490FD8",x"3FC90FD8",x"40490FDC",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"437F0000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"4E6E6B28",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"028000EC",x"02A000C8",x"06C00001",x"0220000B",x"02400000",x"03DC0004",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0004",x"0048A000",x"C4240000",x"06880004",x"86C80650",x"028000C4",x"02A001E0",x"02200001",x"0240FFFF",x"03DC0004",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0004",x"0048A000",x"C4240000",x"06880004",x"86C80684",x"02200001",x"0240FFFF",x"03DC0004",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0004",x"00420000",x"02200001",x"03DC0004",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0004",x"C42002A8",x"02A00368",x"02200003",x"02400000",x"03DC0004",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0004",x"C42A0000",x"0220003C",x"03DC0004",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0004",x"C42A0004",x"028002CC",x"02A00370",x"02200002",x"03DC0004",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0004",x"00E20000",x"02200003",x"02400000",x"03DC0004",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0004",x"C4E20004",x"0048A000",x"C4240000",x"06880004",x"86C80734",x"C1FDFFFC",x"E0200000",x"C1FDFFFC",x"E2200000",x"C1FDFFFC",x"E0200000",x"E0400000",x"E0600000",x"E0800000",x"22221820",x"22441020",x"22660820",x"00224000",x"00226000",x"00228000",x"C1FDFFFC",x"E0200000",x"E0400000",x"E0600000",x"E0800000",x"22221820",x"22441020",x"22660820",x"00224000",x"00226000",x"00228000",x"C43C0004",x"C83C0004",x"C1FDFFFC",x"CC3C0004",x"C03C0004",x"228218A0",x"226210A0",x"224208A0",x"E2800000",x"E2600000",x"E2400000",x"E2200000",x"C1FDFFFC",x"007A0000",x"82200834",x"C45A0000",x"06220001",x"03BA0004",x"82000820",x"00260000",x"C1FDFFFC",x"50220000",x"C1FDFFFC",x"60220000",x"C1FDFFFC",x"C84000C0",x"C86000BC",x"C88000B8",x"C43C0000",x"8E240A10",x"44224000",x"04402000",x"C45C0004",x"8E240898",x"44224000",x"04604000",x"C17DFFFC",x"00260000",x"03DC0010",x"037E000C",x"C57DFFFC",x"8200084C",x"07DC0010",x"820009F8",x"8E26094C",x"8E8208F8",x"C84000B4",x"48442000",x"48442000",x"48442000",x"44424000",x"C86000B0",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"40446000",x"C86000AC",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48262000",x"44242000",x"82000948",x"44262000",x"C84000A8",x"C86000A4",x"48662000",x"48662000",x"44446000",x"C86000A0",x"48662000",x"48662000",x"48662000",x"48662000",x"40446000",x"C860009C",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48262000",x"44242000",x"820009F8",x"8E8209A8",x"C84000B4",x"48442000",x"48442000",x"48442000",x"44424000",x"C86000B0",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"40446000",x"C86000AC",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48262000",x"44242000",x"820009F8",x"44262000",x"C84000A8",x"C86000A4",x"48662000",x"48662000",x"44446000",x"C86000A0",x"48662000",x"48662000",x"48662000",x"48662000",x"40446000",x"C860009C",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48262000",x"44242000",x"02200001",x"C05C0004",x"82420A08",x"82000A0C",x"44202000",x"82000B70",x"8E260AC4",x"8E820A70",x"C84000B4",x"48442000",x"48442000",x"48442000",x"44424000",x"C86000B0",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"40446000",x"C86000AC",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48262000",x"44242000",x"82000AC0",x"44262000",x"C84000A8",x"C86000A4",x"48662000",x"48662000",x"44446000",x"C86000A0",x"48662000",x"48662000",x"48662000",x"48662000",x"40446000",x"C860009C",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48262000",x"44242000",x"82000B70",x"8E820B20",x"C84000B4",x"48442000",x"48442000",x"48442000",x"44424000",x"C86000B0",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"40446000",x"C86000AC",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48262000",x"44242000",x"82000B70",x"44262000",x"C84000A8",x"C86000A4",x"48662000",x"48662000",x"44446000",x"C86000A0",x"48662000",x"48662000",x"48662000",x"48662000",x"40446000",x"C860009C",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48262000",x"44242000",x"02200001",x"C05C0000",x"82420B80",x"C1FDFFFC",x"44202000",x"C1FDFFFC",x"C84000C0",x"C86000BC",x"C88000B8",x"C43C0000",x"8E240D4C",x"44224000",x"04402000",x"C45C0004",x"8E240BD4",x"44224000",x"04604000",x"C17DFFFC",x"00260000",x"03DC0010",x"037E000C",x"C57DFFFC",x"8200084C",x"07DC0010",x"82000D34",x"8E260C88",x"8E820C34",x"C84000B4",x"48442000",x"48442000",x"48442000",x"44424000",x"C86000B0",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"40446000",x"C86000AC",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48262000",x"44242000",x"82000C84",x"44262000",x"C84000A8",x"C86000A4",x"48662000",x"48662000",x"44446000",x"C86000A0",x"48662000",x"48662000",x"48662000",x"48662000",x"40446000",x"C860009C",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48262000",x"44242000",x"82000D34",x"8E820CE4",x"C84000B4",x"48442000",x"48442000",x"48442000",x"44424000",x"C86000B0",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"40446000",x"C86000AC",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48262000",x"44242000",x"82000D34",x"44262000",x"C84000A8",x"C86000A4",x"48662000",x"48662000",x"44446000",x"C86000A0",x"48662000",x"48662000",x"48662000",x"48662000",x"40446000",x"C860009C",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48262000",x"44242000",x"02200001",x"C05C0004",x"82420D44",x"82000D48",x"44202000",x"82000EAC",x"8E260E00",x"8E820DA4",x"C84000A8",x"C86000A4",x"48662000",x"48662000",x"44446000",x"C86000A0",x"48662000",x"48662000",x"48662000",x"48662000",x"40446000",x"C860009C",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48262000",x"44242000",x"82000DFC",x"44262000",x"C84000B4",x"48442000",x"48442000",x"48442000",x"44424000",x"C86000B0",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"40446000",x"C86000AC",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48262000",x"44242000",x"82000EAC",x"8E820E54",x"C84000A8",x"C86000A4",x"48662000",x"48662000",x"44446000",x"C86000A0",x"48662000",x"48662000",x"48662000",x"48662000",x"40446000",x"C860009C",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48262000",x"44242000",x"82000EAC",x"44262000",x"C84000B4",x"48442000",x"48442000",x"48442000",x"44424000",x"C86000B0",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"40446000",x"C86000AC",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48262000",x"44242000",x"02200001",x"C05C0000",x"82420EBC",x"C1FDFFFC",x"44202000",x"C1FDFFFC",x"C8400098",x"8E240F00",x"44224000",x"8E240EDC",x"44224000",x"82000EC4",x"8E020EF8",x"C8600090",x"8E620EF0",x"40224000",x"82000EC4",x"02200001",x"8200084C",x"0220FFFF",x"8200084C",x"8E0210D8",x"C8600090",x"8E620F3C",x"40224000",x"8E240F1C",x"44224000",x"82000EC4",x"8E020F34",x"8E620F2C",x"40224000",x"82000EC4",x"02200001",x"8200084C",x"0220FFFF",x"8200084C",x"C84000C0",x"C86000BC",x"C88000B8",x"8E240F70",x"44224000",x"0220FFFF",x"C17DFFFC",x"03DC0008",x"037E000C",x"C57DFFFC",x"8200084C",x"07DC0008",x"820010D0",x"8E261024",x"8E820FD0",x"C84000B4",x"48442000",x"48442000",x"48442000",x"44424000",x"C86000B0",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"40446000",x"C86000AC",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48262000",x"44242000",x"82001020",x"44262000",x"C84000A8",x"C86000A4",x"48662000",x"48662000",x"44446000",x"C86000A0",x"48662000",x"48662000",x"48662000",x"48662000",x"40446000",x"C860009C",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48262000",x"44242000",x"820010D0",x"8E821080",x"C84000B4",x"48442000",x"48442000",x"48442000",x"44424000",x"C86000B0",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"40446000",x"C86000AC",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48262000",x"44242000",x"820010D0",x"44262000",x"C84000A8",x"C86000A4",x"48662000",x"48662000",x"44446000",x"C86000A0",x"48662000",x"48662000",x"48662000",x"48662000",x"40446000",x"C860009C",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48262000",x"44242000",x"44202000",x"C1FDFFFC",x"C84000C0",x"C86000BC",x"C88000B8",x"8E24110C",x"44224000",x"02200001",x"C17DFFFC",x"03DC0008",x"037E000C",x"C57DFFFC",x"8200084C",x"07DC0008",x"8200126C",x"8E2611C0",x"8E82116C",x"C84000B4",x"48442000",x"48442000",x"48442000",x"44424000",x"C86000B0",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"40446000",x"C86000AC",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48262000",x"44242000",x"820011BC",x"44262000",x"C84000A8",x"C86000A4",x"48662000",x"48662000",x"44446000",x"C86000A0",x"48662000",x"48662000",x"48662000",x"48662000",x"40446000",x"C860009C",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48262000",x"44242000",x"8200126C",x"8E82121C",x"C84000B4",x"48442000",x"48442000",x"48442000",x"44424000",x"C86000B0",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"40446000",x"C86000AC",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48262000",x"44242000",x"8200126C",x"44262000",x"C84000A8",x"C86000A4",x"48662000",x"48662000",x"44446000",x"C86000A0",x"48662000",x"48662000",x"48662000",x"48662000",x"40446000",x"C860009C",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48262000",x"44242000",x"C1FDFFFC",x"C8400098",x"8E2412AC",x"44224000",x"8E241288",x"44224000",x"82001270",x"8E0212A4",x"C8600090",x"8E62129C",x"40224000",x"82001270",x"02200001",x"82000B88",x"0220FFFF",x"82000B88",x"8E021484",x"C8600090",x"8E6212E8",x"40224000",x"8E2412C8",x"44224000",x"82001270",x"8E0212E0",x"8E6212D8",x"40224000",x"82001270",x"02200001",x"82000B88",x"0220FFFF",x"82000B88",x"C84000C0",x"C86000BC",x"C88000B8",x"8E24131C",x"44224000",x"0220FFFF",x"C17DFFFC",x"03DC0008",x"037E000C",x"C57DFFFC",x"8200084C",x"07DC0008",x"8200147C",x"8E2613D0",x"8E821374",x"C84000A8",x"C86000A4",x"48662000",x"48662000",x"44446000",x"C86000A0",x"48662000",x"48662000",x"48662000",x"48662000",x"40446000",x"C860009C",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48262000",x"44242000",x"820013CC",x"44262000",x"C84000B4",x"48442000",x"48442000",x"48442000",x"44424000",x"C86000B0",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"40446000",x"C86000AC",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48262000",x"44242000",x"8200147C",x"8E821424",x"C84000A8",x"C86000A4",x"48662000",x"48662000",x"44446000",x"C86000A0",x"48662000",x"48662000",x"48662000",x"48662000",x"40446000",x"C860009C",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48262000",x"44242000",x"8200147C",x"44262000",x"C84000B4",x"48442000",x"48442000",x"48442000",x"44424000",x"C86000B0",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"40446000",x"C86000AC",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48262000",x"44242000",x"44202000",x"C1FDFFFC",x"C84000C0",x"C86000BC",x"C88000B8",x"8E2414B8",x"44224000",x"02200001",x"C17DFFFC",x"03DC0008",x"037E000C",x"C57DFFFC",x"8200084C",x"07DC0008",x"82001618",x"8E26156C",x"8E821510",x"C84000A8",x"C86000A4",x"48662000",x"48662000",x"44446000",x"C86000A0",x"48662000",x"48662000",x"48662000",x"48662000",x"40446000",x"C860009C",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48262000",x"44242000",x"82001568",x"44262000",x"C84000B4",x"48442000",x"48442000",x"48442000",x"44424000",x"C86000B0",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"40446000",x"C86000AC",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48262000",x"44242000",x"82001618",x"8E8215C0",x"C84000A8",x"C86000A4",x"48662000",x"48662000",x"44446000",x"C86000A0",x"48662000",x"48662000",x"48662000",x"48662000",x"40446000",x"C860009C",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48262000",x"44242000",x"82001618",x"44262000",x"C84000B4",x"48442000",x"48442000",x"48442000",x"44424000",x"C86000B0",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"40446000",x"C86000AC",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48662000",x"48262000",x"44242000",x"C1FDFFFC",x"C8220000",x"48222000",x"C8420004",x"48444000",x"40224000",x"C8420008",x"48444000",x"40224000",x"C43C0000",x"C45C0004",x"C17DFFFC",x"03DC0010",x"037E000C",x"C57DFFFC",x"8200083C",x"07DC0010",x"8A2016A4",x"C03C0004",x"82201688",x"C17DFFFC",x"03DC0010",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0010",x"44202000",x"820016A0",x"C17DFFFC",x"03DC0010",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0010",x"820016A8",x"C82000A8",x"C03C0000",x"C8420000",x"48442000",x"CC420000",x"C8420004",x"48442000",x"CC420004",x"C8420008",x"48242000",x"CC220008",x"C1FDFFFC",x"022001B8",x"C43C0000",x"C17DFFFC",x"03DC000C",x"037E000C",x"C57DFFFC",x"820007C0",x"07DC000C",x"C03C0000",x"CC220000",x"C17DFFFC",x"03DC000C",x"037E000C",x"C57DFFFC",x"820007C0",x"07DC000C",x"C03C0000",x"CC220004",x"C17DFFFC",x"03DC000C",x"037E000C",x"C57DFFFC",x"820007C0",x"07DC000C",x"C03C0000",x"CC220008",x"C17DFFFC",x"03DC000C",x"037E000C",x"C57DFFFC",x"820007C0",x"07DC000C",x"C840008C",x"48224000",x"C8600098",x"CC5C0008",x"CC7C0010",x"CC3C0018",x"8E261794",x"44826000",x"C17DFFFC",x"40208000",x"03DC0028",x"037E000C",x"C57DFFFC",x"82001270",x"07DC0028",x"82001800",x"8E0217E4",x"C8800090",x"8E8217C4",x"40826000",x"C17DFFFC",x"40208000",x"03DC0028",x"037E000C",x"C57DFFFC",x"82001270",x"07DC0028",x"820017E0",x"02200001",x"C17DFFFC",x"03DC0028",x"037E000C",x"C57DFFFC",x"82000B88",x"07DC0028",x"82001800",x"0220FFFF",x"C17DFFFC",x"03DC0028",x"037E000C",x"C57DFFFC",x"82000B88",x"07DC0028",x"C85C0010",x"C87C0018",x"CC3C0020",x"8E641834",x"44664000",x"C17DFFFC",x"40206000",x"03DC0030",x"037E000C",x"C57DFFFC",x"82000EC4",x"07DC0030",x"820018A8",x"8E061888",x"C8800090",x"8E861864",x"40664000",x"C17DFFFC",x"40206000",x"03DC0030",x"037E000C",x"C57DFFFC",x"82000EC4",x"07DC0030",x"82001884",x"02200001",x"C17DFFFC",x"40206000",x"03DC0030",x"037E000C",x"C57DFFFC",x"8200084C",x"07DC0030",x"820018A8",x"0220FFFF",x"C17DFFFC",x"40206000",x"03DC0030",x"037E000C",x"C57DFFFC",x"8200084C",x"07DC0030",x"CC3C0028",x"C17DFFFC",x"03DC0038",x"037E000C",x"C57DFFFC",x"820007C0",x"07DC0038",x"C85C0008",x"48224000",x"C85C0010",x"CC3C0030",x"8E2418FC",x"44624000",x"C17DFFFC",x"40206000",x"03DC0040",x"037E000C",x"C57DFFFC",x"82001270",x"07DC0040",x"82001968",x"8E02194C",x"C8600090",x"8E62192C",x"40624000",x"C17DFFFC",x"40206000",x"03DC0040",x"037E000C",x"C57DFFFC",x"82001270",x"07DC0040",x"82001948",x"02200001",x"C17DFFFC",x"03DC0040",x"037E000C",x"C57DFFFC",x"82000B88",x"07DC0040",x"82001968",x"0220FFFF",x"C17DFFFC",x"03DC0040",x"037E000C",x"C57DFFFC",x"82000B88",x"07DC0040",x"C85C0010",x"C87C0030",x"CC3C0038",x"8E64199C",x"44464000",x"C17DFFFC",x"40204000",x"03DC0048",x"037E000C",x"C57DFFFC",x"82000EC4",x"07DC0048",x"82001A10",x"8E0619F0",x"C8800090",x"8E8619CC",x"40464000",x"C17DFFFC",x"40204000",x"03DC0048",x"037E000C",x"C57DFFFC",x"82000EC4",x"07DC0048",x"820019EC",x"02200001",x"C17DFFFC",x"40206000",x"03DC0048",x"037E000C",x"C57DFFFC",x"8200084C",x"07DC0048",x"82001A10",x"0220FFFF",x"C17DFFFC",x"40206000",x"03DC0048",x"037E000C",x"C57DFFFC",x"8200084C",x"07DC0048",x"0220033C",x"C85C0020",x"48642000",x"C8800088",x"48668000",x"CC620000",x"C8600084",x"C8BC0028",x"486A6000",x"CC620004",x"C87C0038",x"48C46000",x"488C8000",x"CC820008",x"02400324",x"CC640000",x"CC040004",x"44802000",x"CC840008",x"02400330",x"4480A000",x"48282000",x"CC240000",x"44204000",x"CC240004",x"48286000",x"CC240008",x"024001C4",x"C07C0000",x"C8260000",x"C8420000",x"44224000",x"CC240000",x"C8260004",x"C8420004",x"44224000",x"CC240004",x"C8260008",x"C8420008",x"44224000",x"CC240008",x"C1FDFFFC",x"C17DFFFC",x"03DC0008",x"037E000C",x"C57DFFFC",x"82000794",x"07DC0008",x"C17DFFFC",x"03DC0008",x"037E000C",x"C57DFFFC",x"820007C0",x"07DC0008",x"C840008C",x"48224000",x"C8600098",x"CC7C0000",x"CC3C0008",x"CC5C0010",x"8E261B28",x"44826000",x"C17DFFFC",x"40208000",x"03DC0020",x"037E000C",x"C57DFFFC",x"82000EC4",x"07DC0020",x"82001B94",x"8E021B78",x"C8800090",x"8E821B58",x"40826000",x"C17DFFFC",x"40208000",x"03DC0020",x"037E000C",x"C57DFFFC",x"82000EC4",x"07DC0020",x"82001B74",x"02200001",x"C17DFFFC",x"03DC0020",x"037E000C",x"C57DFFFC",x"8200084C",x"07DC0020",x"82001B94",x"0220FFFF",x"C17DFFFC",x"03DC0020",x"037E000C",x"C57DFFFC",x"8200084C",x"07DC0020",x"022001D0",x"44202000",x"CC220004",x"C43C0018",x"C17DFFFC",x"03DC0024",x"037E000C",x"C57DFFFC",x"820007C0",x"07DC0024",x"C85C0010",x"48224000",x"C85C0000",x"C87C0008",x"CC3C0020",x"8E641BF8",x"44664000",x"C17DFFFC",x"40206000",x"03DC0030",x"037E000C",x"C57DFFFC",x"82001270",x"07DC0030",x"82001C6C",x"8E061C4C",x"C8800090",x"8E861C28",x"40664000",x"C17DFFFC",x"40206000",x"03DC0030",x"037E000C",x"C57DFFFC",x"82001270",x"07DC0030",x"82001C48",x"02200001",x"C17DFFFC",x"40206000",x"03DC0030",x"037E000C",x"C57DFFFC",x"82000B88",x"07DC0030",x"82001C6C",x"0220FFFF",x"C17DFFFC",x"40206000",x"03DC0030",x"037E000C",x"C57DFFFC",x"82000B88",x"07DC0030",x"C85C0000",x"C87C0020",x"CC3C0028",x"8E641CA0",x"44864000",x"C17DFFFC",x"40208000",x"03DC0038",x"037E000C",x"C57DFFFC",x"82000EC4",x"07DC0038",x"82001D14",x"8E061CF4",x"C8800090",x"8E861CD0",x"40864000",x"C17DFFFC",x"40208000",x"03DC0038",x"037E000C",x"C57DFFFC",x"82000EC4",x"07DC0038",x"82001CF0",x"02200001",x"C17DFFFC",x"40206000",x"03DC0038",x"037E000C",x"C57DFFFC",x"8200084C",x"07DC0038",x"82001D14",x"0220FFFF",x"C17DFFFC",x"40206000",x"03DC0038",x"037E000C",x"C57DFFFC",x"8200084C",x"07DC0038",x"C85C0028",x"48242000",x"C03C0018",x"CC220000",x"C83C0000",x"C87C0020",x"8E621D50",x"44262000",x"C17DFFFC",x"03DC0038",x"037E000C",x"C57DFFFC",x"82001270",x"07DC0038",x"82001DC8",x"8E061DA4",x"C8800090",x"8E861D7C",x"40262000",x"C17DFFFC",x"03DC0038",x"037E000C",x"C57DFFFC",x"82001270",x"07DC0038",x"82001DA0",x"02400001",x"C17DFFFC",x"00240000",x"40206000",x"03DC0038",x"037E000C",x"C57DFFFC",x"82000B88",x"07DC0038",x"82001DC8",x"0240FFFF",x"C17DFFFC",x"00240000",x"40206000",x"03DC0038",x"037E000C",x"C57DFFFC",x"82000B88",x"07DC0038",x"C85C0028",x"48242000",x"C03C0018",x"CC220008",x"022001DC",x"C43C0030",x"C17DFFFC",x"03DC003C",x"037E000C",x"C57DFFFC",x"820007C0",x"07DC003C",x"C03C0030",x"CC220000",x"C1FDFFFC",x"C8240000",x"C8400098",x"C43C0000",x"CC5C0008",x"C45C0010",x"8E241E3C",x"44224000",x"C17DFFFC",x"03DC001C",x"037E000C",x"C57DFFFC",x"82001270",x"07DC001C",x"82001EAC",x"8E021E8C",x"C8600090",x"8E621E68",x"40224000",x"C17DFFFC",x"03DC001C",x"037E000C",x"C57DFFFC",x"82001270",x"07DC001C",x"82001E88",x"02600001",x"C17DFFFC",x"00260000",x"03DC001C",x"037E000C",x"C57DFFFC",x"82000B88",x"07DC001C",x"82001EAC",x"0260FFFF",x"C17DFFFC",x"00260000",x"03DC001C",x"037E000C",x"C57DFFFC",x"82000B88",x"07DC001C",x"C03C0010",x"C8420000",x"C87C0008",x"CC3C0018",x"8E461EE4",x"44446000",x"C17DFFFC",x"40204000",x"03DC0028",x"037E000C",x"C57DFFFC",x"82000EC4",x"07DC0028",x"82001F60",x"8E041F3C",x"C8800090",x"8E841F14",x"40446000",x"C17DFFFC",x"40204000",x"03DC0028",x"037E000C",x"C57DFFFC",x"82000EC4",x"07DC0028",x"82001F38",x"02400001",x"C17DFFFC",x"00240000",x"40204000",x"03DC0028",x"037E000C",x"C57DFFFC",x"8200084C",x"07DC0028",x"82001F60",x"0240FFFF",x"C17DFFFC",x"00240000",x"40204000",x"03DC0028",x"037E000C",x"C57DFFFC",x"8200084C",x"07DC0028",x"C03C0010",x"C8420004",x"C87C0008",x"CC3C0020",x"8E461F98",x"44446000",x"C17DFFFC",x"40204000",x"03DC0030",x"037E000C",x"C57DFFFC",x"82001270",x"07DC0030",x"82002014",x"8E041FF0",x"C8800090",x"8E841FC8",x"40446000",x"C17DFFFC",x"40204000",x"03DC0030",x"037E000C",x"C57DFFFC",x"82001270",x"07DC0030",x"82001FEC",x"02400001",x"C17DFFFC",x"00240000",x"40204000",x"03DC0030",x"037E000C",x"C57DFFFC",x"82000B88",x"07DC0030",x"82002014",x"0240FFFF",x"C17DFFFC",x"00240000",x"40204000",x"03DC0030",x"037E000C",x"C57DFFFC",x"82000B88",x"07DC0030",x"C03C0010",x"C8420004",x"C87C0008",x"CC3C0028",x"8E46204C",x"44446000",x"C17DFFFC",x"40204000",x"03DC0038",x"037E000C",x"C57DFFFC",x"82000EC4",x"07DC0038",x"820020C8",x"8E0420A4",x"C8800090",x"8E84207C",x"40446000",x"C17DFFFC",x"40204000",x"03DC0038",x"037E000C",x"C57DFFFC",x"82000EC4",x"07DC0038",x"820020A0",x"02400001",x"C17DFFFC",x"00240000",x"40204000",x"03DC0038",x"037E000C",x"C57DFFFC",x"8200084C",x"07DC0038",x"820020C8",x"0240FFFF",x"C17DFFFC",x"00240000",x"40204000",x"03DC0038",x"037E000C",x"C57DFFFC",x"8200084C",x"07DC0038",x"C03C0010",x"C8420008",x"C87C0008",x"CC3C0030",x"8E462100",x"44446000",x"C17DFFFC",x"40204000",x"03DC0040",x"037E000C",x"C57DFFFC",x"82001270",x"07DC0040",x"8200217C",x"8E042158",x"C8800090",x"8E842130",x"40446000",x"C17DFFFC",x"40204000",x"03DC0040",x"037E000C",x"C57DFFFC",x"82001270",x"07DC0040",x"82002154",x"02400001",x"C17DFFFC",x"00240000",x"40204000",x"03DC0040",x"037E000C",x"C57DFFFC",x"82000B88",x"07DC0040",x"8200217C",x"0240FFFF",x"C17DFFFC",x"00240000",x"40204000",x"03DC0040",x"037E000C",x"C57DFFFC",x"82000B88",x"07DC0040",x"C03C0010",x"C8420008",x"C87C0008",x"CC3C0038",x"8E4621B4",x"44446000",x"C17DFFFC",x"40204000",x"03DC0048",x"037E000C",x"C57DFFFC",x"82000EC4",x"07DC0048",x"82002230",x"8E04220C",x"C8800090",x"8E8421E4",x"40446000",x"C17DFFFC",x"40204000",x"03DC0048",x"037E000C",x"C57DFFFC",x"82000EC4",x"07DC0048",x"82002208",x"02400001",x"C17DFFFC",x"00240000",x"40204000",x"03DC0048",x"037E000C",x"C57DFFFC",x"8200084C",x"07DC0048",x"82002230",x"0240FFFF",x"C17DFFFC",x"00240000",x"40204000",x"03DC0048",x"037E000C",x"C57DFFFC",x"8200084C",x"07DC0048",x"C85C0038",x"C87C0028",x"48864000",x"C8BC0030",x"C8DC0020",x"48ECA000",x"490E4000",x"C93C0018",x"49522000",x"45114000",x"4952A000",x"49744000",x"498C2000",x"41778000",x"49862000",x"48EE2000",x"49B24000",x"40EFA000",x"48342000",x"484C4000",x"44224000",x"4440A000",x"48AC6000",x"48726000",x"C03C0000",x"C8C20000",x"C9220004",x"C9420008",x"49A88000",x"49ADA000",x"49D98000",x"49D3C000",x"41BBC000",x"49C44000",x"49D5C000",x"41BBC000",x"CDA20000",x"49B10000",x"49ADA000",x"49CEE000",x"49D3C000",x"41BBC000",x"49CAA000",x"49D5C000",x"41BBC000",x"CDA20004",x"49B76000",x"49ADA000",x"49C22000",x"49D3C000",x"41BBC000",x"49C66000",x"49D5C000",x"41BBC000",x"CDA20008",x"C9A00080",x"49CD0000",x"49DD6000",x"49F2E000",x"49FE2000",x"41DDE000",x"49F4A000",x"49FE6000",x"41DDE000",x"49DBC000",x"C03C0010",x"CDC20000",x"488C8000",x"48C96000",x"49338000",x"48322000",x"402C2000",x"48544000",x"48646000",x"40226000",x"483A2000",x"CC220004",x"48290000",x"4872E000",x"40226000",x"4844A000",x"40224000",x"483A2000",x"CC220008",x"C1FDFFFC",x"C43C0000",x"C17DFFFC",x"03DC000C",x"037E000C",x"C57DFFFC",x"82000794",x"07DC000C",x"0240FFFF",x"82242928",x"C43C0004",x"C17DFFFC",x"03DC0010",x"037E000C",x"C57DFFFC",x"82000794",x"07DC0010",x"C43C0008",x"C17DFFFC",x"03DC0014",x"037E000C",x"C57DFFFC",x"82000794",x"07DC0014",x"C43C000C",x"C17DFFFC",x"03DC0018",x"037E000C",x"C57DFFFC",x"82000794",x"07DC0018",x"02400003",x"40200000",x"C43C0010",x"CC3C0018",x"C17DFFFC",x"00240000",x"03DC0028",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0028",x"C43C0020",x"C17DFFFC",x"03DC002C",x"037E000C",x"C57DFFFC",x"820007C0",x"07DC002C",x"C03C0020",x"CC220000",x"C17DFFFC",x"03DC002C",x"037E000C",x"C57DFFFC",x"820007C0",x"07DC002C",x"C03C0020",x"CC220004",x"C17DFFFC",x"03DC002C",x"037E000C",x"C57DFFFC",x"820007C0",x"07DC002C",x"C03C0020",x"CC220008",x"02400003",x"C83C0018",x"C17DFFFC",x"00240000",x"03DC002C",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC002C",x"C43C0024",x"C17DFFFC",x"03DC0030",x"037E000C",x"C57DFFFC",x"820007C0",x"07DC0030",x"C03C0024",x"CC220000",x"C17DFFFC",x"03DC0030",x"037E000C",x"C57DFFFC",x"820007C0",x"07DC0030",x"C03C0024",x"CC220004",x"C17DFFFC",x"03DC0030",x"037E000C",x"C57DFFFC",x"820007C0",x"07DC0030",x"C03C0024",x"CC220008",x"C17DFFFC",x"03DC0030",x"037E000C",x"C57DFFFC",x"820007C0",x"07DC0030",x"8E202538",x"02200000",x"8200253C",x"02200001",x"02400002",x"C85C0018",x"CC3C0028",x"C43C0030",x"C17DFFFC",x"00240000",x"40204000",x"03DC003C",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC003C",x"C43C0034",x"C17DFFFC",x"03DC0040",x"037E000C",x"C57DFFFC",x"820007C0",x"07DC0040",x"C03C0034",x"CC220000",x"C17DFFFC",x"03DC0040",x"037E000C",x"C57DFFFC",x"820007C0",x"07DC0040",x"C03C0034",x"CC220004",x"02400003",x"C83C0018",x"C17DFFFC",x"00240000",x"03DC0040",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0040",x"C43C0038",x"C17DFFFC",x"03DC0044",x"037E000C",x"C57DFFFC",x"820007C0",x"07DC0044",x"C03C0038",x"CC220000",x"C17DFFFC",x"03DC0044",x"037E000C",x"C57DFFFC",x"820007C0",x"07DC0044",x"C03C0038",x"CC220004",x"C17DFFFC",x"03DC0044",x"037E000C",x"C57DFFFC",x"820007C0",x"07DC0044",x"C03C0038",x"CC220008",x"02400003",x"C83C0018",x"C17DFFFC",x"00240000",x"03DC0044",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0044",x"C05C0010",x"824026E8",x"C43C003C",x"C17DFFFC",x"03DC0048",x"037E000C",x"C57DFFFC",x"820007C0",x"07DC0048",x"C840008C",x"48224000",x"C03C003C",x"CC220000",x"CC5C0040",x"C17DFFFC",x"03DC0050",x"037E000C",x"C57DFFFC",x"820007C0",x"07DC0050",x"C85C0040",x"48224000",x"C03C003C",x"CC220004",x"C17DFFFC",x"03DC0050",x"037E000C",x"C57DFFFC",x"820007C0",x"07DC0050",x"C85C0040",x"48224000",x"C03C003C",x"CC220008",x"820026E8",x"02400002",x"C07C0008",x"826426FC",x"C05C0030",x"82002700",x"02400001",x"02800004",x"C83C0018",x"C45C0048",x"C43C003C",x"C17DFFFC",x"00280000",x"03DC0054",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0054",x"005A0000",x"03BA002C",x"C4240028",x"C03C003C",x"C4240024",x"C07C0038",x"C4640020",x"C07C0034",x"C464001C",x"C07C0048",x"C4640018",x"C07C0024",x"C4640014",x"C07C0020",x"C4640010",x"C09C0010",x"C484000C",x"C0BC000C",x"C4A40008",x"C0BC0008",x"C4A40004",x"C0DC0004",x"C4C40000",x"02C000C8",x"C0FC0000",x"22EE0220",x"D44CE000",x"02400003",x"82A427E0",x"02400002",x"82A427AC",x"820027DC",x"C83C0028",x"8E2027BC",x"02400001",x"820027C0",x"02400000",x"C17DFFFC",x"00260000",x"03DC0054",x"037E000C",x"C57DFFFC",x"8200161C",x"07DC0054",x"820028F4",x"C8260000",x"8A202830",x"8A202800",x"8E0227F8",x"C840007C",x"820027FC",x"C84000A8",x"82002804",x"40400000",x"48222000",x"CC5C0050",x"C17DFFFC",x"03DC0060",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0060",x"C85C0050",x"48242000",x"82002834",x"40200000",x"C03C0020",x"CC220000",x"C8220004",x"8A20288C",x"8A20285C",x"8E022854",x"C840007C",x"82002858",x"C84000A8",x"82002860",x"40400000",x"48222000",x"CC5C0058",x"C17DFFFC",x"03DC0068",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0068",x"C85C0058",x"48242000",x"82002890",x"40200000",x"C03C0020",x"CC220004",x"C8220008",x"8A2028E8",x"8A2028B8",x"8E0228B0",x"C840007C",x"820028B4",x"C84000A8",x"820028BC",x"40400000",x"48222000",x"CC5C0060",x"C17DFFFC",x"03DC0070",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0070",x"C85C0060",x"48242000",x"820028EC",x"40200000",x"C03C0020",x"CC220008",x"C03C0010",x"82202920",x"C03C0020",x"C05C003C",x"C17DFFFC",x"03DC0070",x"037E000C",x"C57DFFFC",x"82001E04",x"07DC0070",x"82002920",x"02200001",x"C1FDFFFC",x"02200000",x"C1FDFFFC",x"0240003C",x"8624293C",x"C1FDFFFC",x"C43C0000",x"C17DFFFC",x"03DC000C",x"037E000C",x"C57DFFFC",x"82002384",x"07DC000C",x"82202A34",x"C03C0000",x"02220001",x"0240003C",x"86242970",x"C1FDFFFC",x"C43C0004",x"C17DFFFC",x"03DC0010",x"037E000C",x"C57DFFFC",x"82002384",x"07DC0010",x"82202A24",x"C03C0004",x"02220001",x"0240003C",x"862429A4",x"C1FDFFFC",x"C43C0008",x"C17DFFFC",x"03DC0014",x"037E000C",x"C57DFFFC",x"82002384",x"07DC0014",x"82202A14",x"C03C0008",x"02220001",x"0240003C",x"862429D8",x"C1FDFFFC",x"C43C000C",x"C17DFFFC",x"03DC0018",x"037E000C",x"C57DFFFC",x"82002384",x"07DC0018",x"82202A04",x"C03C000C",x"02220001",x"82002930",x"022000C4",x"C05C000C",x"C4420000",x"C1FDFFFC",x"022000C4",x"C05C0008",x"C4420000",x"C1FDFFFC",x"022000C4",x"C05C0004",x"C4420000",x"C1FDFFFC",x"022000C4",x"C05C0000",x"C4420000",x"C1FDFFFC",x"C43C0000",x"C17DFFFC",x"03DC000C",x"037E000C",x"C57DFFFC",x"82000794",x"07DC000C",x"0240FFFF",x"82242BDC",x"C05C0000",x"02640001",x"C43C0004",x"C47C0008",x"C17DFFFC",x"03DC0014",x"037E000C",x"C57DFFFC",x"82000794",x"07DC0014",x"0240FFFF",x"82242BA4",x"C05C0008",x"02640001",x"C43C000C",x"C47C0010",x"C17DFFFC",x"03DC001C",x"037E000C",x"C57DFFFC",x"82000794",x"07DC001C",x"0240FFFF",x"82242B6C",x"C05C0010",x"02640001",x"C43C0014",x"C47C0018",x"C17DFFFC",x"03DC0024",x"037E000C",x"C57DFFFC",x"82000794",x"07DC0024",x"0240FFFF",x"82242B34",x"C05C0018",x"02640001",x"C43C001C",x"C17DFFFC",x"00260000",x"03DC0028",x"037E000C",x"C57DFFFC",x"82002A44",x"07DC0028",x"C05C0018",x"22440220",x"C07C001C",x"D4624000",x"82002B58",x"C03C0018",x"02220001",x"0240FFFF",x"C17DFFFC",x"03DC0028",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0028",x"C05C0010",x"22440220",x"C07C0014",x"D4624000",x"82002B90",x"C03C0010",x"02220001",x"0240FFFF",x"C17DFFFC",x"03DC0028",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0028",x"C05C0008",x"22440220",x"C07C000C",x"D4624000",x"82002BC8",x"C03C0008",x"02220001",x"0240FFFF",x"C17DFFFC",x"03DC0028",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0028",x"C05C0000",x"22440220",x"C07C0004",x"D4624000",x"C1FDFFFC",x"C03C0000",x"02220001",x"0240FFFF",x"8200081C",x"C43C0000",x"C17DFFFC",x"03DC000C",x"037E000C",x"C57DFFFC",x"82000794",x"07DC000C",x"0240FFFF",x"82242CE4",x"C43C0004",x"C17DFFFC",x"03DC0010",x"037E000C",x"C57DFFFC",x"82000794",x"07DC0010",x"0240FFFF",x"82242CB4",x"C43C0008",x"C17DFFFC",x"03DC0014",x"037E000C",x"C57DFFFC",x"82000794",x"07DC0014",x"0240FFFF",x"82242C88",x"02400003",x"C43C000C",x"C17DFFFC",x"00240000",x"03DC0018",x"037E000C",x"C57DFFFC",x"82002A44",x"07DC0018",x"C05C000C",x"C4420008",x"82002CA8",x"02200003",x"0240FFFF",x"C17DFFFC",x"03DC0018",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0018",x"C05C0008",x"C4420004",x"82002CD4",x"02200002",x"0240FFFF",x"C17DFFFC",x"03DC0018",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0018",x"C05C0004",x"C4420000",x"00420000",x"82002D08",x"02200001",x"0240FFFF",x"C17DFFFC",x"03DC0018",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0018",x"00420000",x"C0240000",x"0260FFFF",x"82262E68",x"C03C0000",x"02620001",x"C45C0010",x"C47C0014",x"C17DFFFC",x"03DC0020",x"037E000C",x"C57DFFFC",x"82000794",x"07DC0020",x"0240FFFF",x"82242DC8",x"C43C0018",x"C17DFFFC",x"03DC0024",x"037E000C",x"C57DFFFC",x"82000794",x"07DC0024",x"0240FFFF",x"82242D98",x"02400002",x"C43C001C",x"C17DFFFC",x"00240000",x"03DC0028",x"037E000C",x"C57DFFFC",x"82002A44",x"07DC0028",x"C05C001C",x"C4420004",x"82002DB8",x"02200002",x"0240FFFF",x"C17DFFFC",x"03DC0028",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0028",x"C05C0018",x"C4420000",x"00420000",x"82002DEC",x"02200001",x"0240FFFF",x"C17DFFFC",x"03DC0028",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0028",x"00420000",x"C0240000",x"0260FFFF",x"82262E34",x"C03C0014",x"02620001",x"C45C0020",x"C17DFFFC",x"00260000",x"03DC002C",x"037E000C",x"C57DFFFC",x"82002BEC",x"07DC002C",x"C05C0014",x"22440220",x"C07C0020",x"D4624000",x"82002E54",x"C03C0014",x"02220001",x"C17DFFFC",x"03DC002C",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC002C",x"C05C0000",x"22440220",x"C07C0010",x"D4624000",x"C1FDFFFC",x"C03C0000",x"02220001",x"8200081C",x"C43C0000",x"C17DFFFC",x"03DC000C",x"037E000C",x"C57DFFFC",x"82000794",x"07DC000C",x"0240FFFF",x"82242F68",x"C43C0004",x"C17DFFFC",x"03DC0010",x"037E000C",x"C57DFFFC",x"82000794",x"07DC0010",x"0240FFFF",x"82242F3C",x"C43C0008",x"C17DFFFC",x"03DC0014",x"037E000C",x"C57DFFFC",x"82000794",x"07DC0014",x"0240FFFF",x"82242F10",x"02400003",x"C43C000C",x"C17DFFFC",x"00240000",x"03DC0018",x"037E000C",x"C57DFFFC",x"82002A44",x"07DC0018",x"C05C000C",x"C4420008",x"82002F30",x"02200003",x"0240FFFF",x"C17DFFFC",x"03DC0018",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0018",x"C05C0008",x"C4420004",x"82002F5C",x"02200002",x"0240FFFF",x"C17DFFFC",x"03DC0018",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0018",x"C05C0004",x"C4420000",x"82002F88",x"02200001",x"0240FFFF",x"C17DFFFC",x"03DC0018",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0018",x"C0420000",x"0260FFFF",x"82463178",x"024001E0",x"C07C0000",x"22860220",x"D4248000",x"02260001",x"C45C0010",x"C43C0014",x"C17DFFFC",x"03DC0020",x"037E000C",x"C57DFFFC",x"82000794",x"07DC0020",x"0240FFFF",x"82243050",x"C43C0018",x"C17DFFFC",x"03DC0024",x"037E000C",x"C57DFFFC",x"82000794",x"07DC0024",x"0240FFFF",x"82243024",x"02400002",x"C43C001C",x"C17DFFFC",x"00240000",x"03DC0028",x"037E000C",x"C57DFFFC",x"82002A44",x"07DC0028",x"C05C001C",x"C4420004",x"82003044",x"02200002",x"0240FFFF",x"C17DFFFC",x"03DC0028",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0028",x"C05C0018",x"C4420000",x"82003070",x"02200001",x"0240FFFF",x"C17DFFFC",x"03DC0028",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0028",x"C0420000",x"0260FFFF",x"82463174",x"C05C0014",x"22640220",x"C09C0010",x"D4286000",x"02240001",x"C43C0020",x"C17DFFFC",x"03DC002C",x"037E000C",x"C57DFFFC",x"82000794",x"07DC002C",x"0240FFFF",x"822430E4",x"02400001",x"C43C0024",x"C17DFFFC",x"00240000",x"03DC0030",x"037E000C",x"C57DFFFC",x"82002A44",x"07DC0030",x"C05C0024",x"C4420000",x"82003104",x"02200001",x"0240FFFF",x"C17DFFFC",x"03DC0030",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0030",x"C0420000",x"0260FFFF",x"82463170",x"C05C0020",x"22640220",x"C09C0010",x"D4286000",x"02240001",x"02400000",x"C43C0028",x"C17DFFFC",x"00240000",x"03DC0034",x"037E000C",x"C57DFFFC",x"82002A44",x"07DC0034",x"C0420000",x"0260FFFF",x"8246316C",x"C05C0028",x"22640220",x"C09C0010",x"D4286000",x"02240001",x"82002E74",x"C1FDFFFC",x"C1FDFFFC",x"C1FDFFFC",x"C1FDFFFC",x"22C60220",x"D884C000",x"8A80329C",x"C0C20010",x"C0220018",x"8E80319C",x"02E00000",x"820031A0",x"02E00001",x"822031B8",x"8E8031B0",x"02200001",x"820031B4",x"02200000",x"820031BC",x"002E0000",x"22660220",x"D8AC6000",x"822031CC",x"820031D0",x"44A0A000",x"442A2000",x"CC7C0000",x"C4BC0008",x"C4DC000C",x"CC5C0010",x"C45C0018",x"C49C001C",x"CC3C0020",x"C17DFFFC",x"40208000",x"03DC0030",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0030",x"C85C0020",x"48242000",x"C03C001C",x"22420220",x"C07C0018",x"D8464000",x"48424000",x"C87C0010",x"40446000",x"8E403238",x"8200323C",x"44404000",x"22220220",x"C05C000C",x"D8642000",x"8E463254",x"02200000",x"C1FDFFFC",x"C03C0008",x"22820220",x"D8468000",x"48424000",x"C87C0000",x"40446000",x"8E403274",x"82003278",x"44404000",x"22220220",x"D8642000",x"8E46328C",x"02200000",x"C1FDFFFC",x"022002AC",x"CC220000",x"02200001",x"C1FDFFFC",x"02200000",x"C1FDFFFC",x"C0220010",x"C8840000",x"C8A20000",x"4888A000",x"C8A40004",x"C8C20004",x"48AAC000",x"4088A000",x"C8A40008",x"C8C20008",x"48AAC000",x"4088A000",x"8E0832E0",x"02200000",x"C1FDFFFC",x"024002AC",x"C8A20000",x"482A2000",x"C8A20004",x"484A4000",x"40224000",x"C8420008",x"48446000",x"40224000",x"44202000",x"C45C0000",x"CC3C0008",x"C17DFFFC",x"40208000",x"03DC0018",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0018",x"C85C0008",x"48242000",x"C03C0000",x"CC220000",x"02200001",x"C1FDFFFC",x"48822000",x"C0420010",x"C8A40000",x"4888A000",x"48A44000",x"C0420010",x"C8C40004",x"48AAC000",x"4088A000",x"48A66000",x"C0420010",x"C8C40008",x"48AAC000",x"4088A000",x"C042000C",x"824033C4",x"48A46000",x"C0420024",x"C8C40000",x"48AAC000",x"4088A000",x"48662000",x"C0420024",x"C8A40004",x"4866A000",x"40686000",x"48224000",x"C0220024",x"C8420008",x"48224000",x"40262000",x"C1FDFFFC",x"40208000",x"C1FDFFFC",x"48E28000",x"C0420010",x"C9040000",x"48EF0000",x"4904A000",x"C0420010",x"C9240004",x"49112000",x"40EF0000",x"4906C000",x"C0420010",x"C9240008",x"49112000",x"40EF0000",x"C042000C",x"82403498",x"4906A000",x"4924C000",x"41112000",x"C0420024",x"C9240000",x"49112000",x"48C2C000",x"48668000",x"406C6000",x"C0420024",x"C8C40004",x"4866C000",x"40706000",x"4822A000",x"48448000",x"40224000",x"C0220024",x"C8420008",x"48224000",x"40262000",x"C8400080",x"CCFC0000",x"CC3C0008",x"C17DFFFC",x"40204000",x"03DC0018",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0018",x"C85C0008",x"48242000",x"C85C0000",x"40242000",x"C1FDFFFC",x"4020E000",x"C1FDFFFC",x"C8840000",x"C8A40004",x"C8C40008",x"48E88000",x"C0620010",x"C9060000",x"48EF0000",x"490AA000",x"C0620010",x"C9260004",x"49112000",x"40EF0000",x"490CC000",x"C0620010",x"C9260008",x"49112000",x"40EF0000",x"C062000C",x"8260352C",x"490AC000",x"C0620024",x"C9260000",x"49112000",x"40EF0000",x"48CC8000",x"C0620024",x"C9060004",x"48CD0000",x"40CEC000",x"4888A000",x"C0620024",x"C8A60008",x"4888A000",x"408C8000",x"82003530",x"4080E000",x"8A8036CC",x"C8A40000",x"C8C40004",x"C8E40008",x"CC9C0000",x"CC7C0008",x"CC5C0010",x"C43C0018",x"CC3C0020",x"C17DFFFC",x"40802000",x"4020A000",x"40A04000",x"4040C000",x"40C06000",x"4060E000",x"03DC0030",x"037E000C",x"C57DFFFC",x"820033CC",x"07DC0030",x"C85C0020",x"48644000",x"C03C0018",x"C0420010",x"C8840000",x"48668000",x"C89C0010",x"48A88000",x"C0420010",x"C8C40004",x"48AAC000",x"4066A000",x"C8BC0008",x"48CAA000",x"C0420010",x"C8E40008",x"48CCE000",x"4066C000",x"C042000C",x"82403614",x"48C8A000",x"C0420024",x"C8E40000",x"48CCE000",x"4066C000",x"48AA4000",x"C0420024",x"C8C40004",x"48AAC000",x"4066A000",x"48448000",x"C0420024",x"C8840008",x"48448000",x"40464000",x"82003618",x"40406000",x"C0420004",x"02600003",x"82463628",x"82003630",x"C86000A8",x"44446000",x"48622000",x"C89C0000",x"48484000",x"44464000",x"8E04364C",x"02200000",x"C1FDFFFC",x"CC3C0028",x"C17DFFFC",x"40204000",x"03DC0038",x"037E000C",x"C57DFFFC",x"8200083C",x"07DC0038",x"C03C0018",x"C0220018",x"8220367C",x"82003680",x"44202000",x"022002AC",x"C85C0028",x"44224000",x"C85C0000",x"C43C0030",x"CC3C0038",x"C17DFFFC",x"40204000",x"03DC0048",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0048",x"C85C0038",x"48242000",x"C03C0030",x"CC220000",x"02200001",x"C1FDFFFC",x"02200000",x"C1FDFFFC",x"028000C8",x"22220220",x"D0282000",x"C8260000",x"C0820014",x"C8480000",x"44224000",x"C8460004",x"C0820014",x"C8680004",x"44446000",x"C8660008",x"C0620014",x"C8860008",x"44668000",x"C0620004",x"02800001",x"826837C8",x"02800002",x"82683728",x"820034A0",x"C0220010",x"C8840000",x"C8A20000",x"4888A000",x"C8A40004",x"C8C20004",x"48AAC000",x"4088A000",x"C8A40008",x"C8C20008",x"48AAC000",x"4088A000",x"8E083764",x"02200000",x"C1FDFFFC",x"024002AC",x"C8A20000",x"482A2000",x"C8A20004",x"484A4000",x"40224000",x"C8420008",x"48446000",x"40224000",x"44202000",x"C45C0000",x"CC3C0008",x"C17DFFFC",x"40208000",x"03DC0018",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0018",x"C85C0008",x"48242000",x"C03C0000",x"CC220000",x"02200001",x"C1FDFFFC",x"02600000",x"02800001",x"02A00002",x"CC3C0010",x"CC7C0018",x"CC5C0020",x"C45C0028",x"C43C002C",x"C17DFFFC",x"03DC0038",x"037E000C",x"C57DFFFC",x"8200317C",x"07DC0038",x"8220380C",x"02200001",x"C1FDFFFC",x"02600001",x"02800002",x"02A00000",x"C83C0020",x"C85C0018",x"C87C0010",x"C03C002C",x"C05C0028",x"C17DFFFC",x"03DC0038",x"037E000C",x"C57DFFFC",x"8200317C",x"07DC0038",x"82203850",x"02200002",x"C1FDFFFC",x"02600002",x"02800000",x"02A00001",x"C83C0018",x"C85C0010",x"C87C0020",x"C03C002C",x"C05C0028",x"C17DFFFC",x"03DC0038",x"037E000C",x"C57DFFFC",x"8200317C",x"07DC0038",x"82203894",x"02200003",x"C1FDFFFC",x"02200000",x"C1FDFFFC",x"C8860000",x"44882000",x"C8A60004",x"4888A000",x"C8A40004",x"48A8A000",x"40AA4000",x"8EA038C0",x"820038C4",x"44A0A000",x"C0820010",x"C8C80004",x"8EAC38D8",x"02800000",x"82003918",x"C8A40008",x"48A8A000",x"40AA6000",x"8EA038EC",x"820038F0",x"44A0A000",x"C0820010",x"C8C80008",x"8EAC3904",x"02800000",x"82003918",x"C8A60004",x"8AA03914",x"02800001",x"82003918",x"02800000",x"8280392C",x"022002AC",x"CC820000",x"02200001",x"C1FDFFFC",x"C8860008",x"44884000",x"C8A6000C",x"4888A000",x"C8A40000",x"48A8A000",x"40AA2000",x"8EA03950",x"82003954",x"44A0A000",x"C0820010",x"C8C80000",x"8EAC3968",x"02800000",x"820039A8",x"C8A40008",x"48A8A000",x"40AA6000",x"8EA0397C",x"82003980",x"44A0A000",x"C0820010",x"C8C80008",x"8EAC3994",x"02800000",x"820039A8",x"C8A6000C",x"8AA039A4",x"02800001",x"820039A8",x"02800000",x"828039BC",x"022002AC",x"CC820000",x"02200002",x"C1FDFFFC",x"C8860010",x"44686000",x"C8860014",x"48668000",x"C8840000",x"48868000",x"40282000",x"8E2039E0",x"820039E4",x"44202000",x"C0820010",x"C8880000",x"8E2839F8",x"02200000",x"82003A38",x"C8240004",x"48262000",x"40224000",x"8E203A0C",x"82003A10",x"44202000",x"C0220010",x"C8420004",x"8E243A24",x"02200000",x"82003A38",x"C8260014",x"8A203A34",x"02200001",x"82003A38",x"02200000",x"82203A4C",x"022002AC",x"CC620000",x"02200003",x"C1FDFFFC",x"02200000",x"C1FDFFFC",x"C8840000",x"8A803BCC",x"C8A40004",x"48AA2000",x"C8C40008",x"48CC4000",x"40AAC000",x"C8C4000C",x"48CC6000",x"40AAC000",x"48C22000",x"C0620010",x"C8E60000",x"48CCE000",x"48E44000",x"C0620010",x"C9060004",x"48EF0000",x"40CCE000",x"48E66000",x"C0620010",x"C9060008",x"48EF0000",x"40CCE000",x"C062000C",x"82603AFC",x"48E46000",x"C0620024",x"C9060000",x"48EF0000",x"40CCE000",x"48662000",x"C0620024",x"C8E60004",x"4866E000",x"406C6000",x"48224000",x"C0620024",x"C8460008",x"48224000",x"40262000",x"82003B00",x"4020C000",x"C0620004",x"02800003",x"82683B10",x"82003B18",x"C84000A8",x"44224000",x"484AA000",x"48282000",x"44242000",x"8E023B30",x"02200000",x"C1FDFFFC",x"C0220018",x"82203B80",x"022002AC",x"C43C0000",x"C45C0004",x"CCBC0008",x"C17DFFFC",x"03DC0018",x"037E000C",x"C57DFFFC",x"8200083C",x"07DC0018",x"C85C0008",x"40242000",x"C03C0004",x"C8420010",x"48224000",x"C03C0000",x"CC220000",x"82003BC4",x"022002AC",x"C43C0010",x"C45C0004",x"CCBC0008",x"C17DFFFC",x"03DC001C",x"037E000C",x"C57DFFFC",x"8200083C",x"07DC001C",x"C85C0008",x"44242000",x"C03C0004",x"C8420010",x"48224000",x"C03C0010",x"CC220000",x"02200001",x"C1FDFFFC",x"02200000",x"C1FDFFFC",x"C8840000",x"8A803CBC",x"C8A40004",x"482A2000",x"C8A40008",x"484A4000",x"40224000",x"C844000C",x"48446000",x"40224000",x"C846000C",x"48622000",x"48484000",x"44464000",x"8E043C18",x"02200000",x"C1FDFFFC",x"C0220018",x"82203C6C",x"022002AC",x"C43C0000",x"C45C0004",x"CC3C0008",x"C17DFFFC",x"40204000",x"03DC0018",x"037E000C",x"C57DFFFC",x"8200083C",x"07DC0018",x"C85C0008",x"40242000",x"C03C0004",x"C8420010",x"48224000",x"C03C0000",x"CC220000",x"82003CB4",x"022002AC",x"C43C0010",x"C45C0004",x"CC3C0008",x"C17DFFFC",x"40204000",x"03DC001C",x"037E000C",x"C57DFFFC",x"8200083C",x"07DC001C",x"C85C0008",x"44242000",x"C03C0004",x"C8420010",x"48224000",x"C03C0010",x"CC220000",x"02200001",x"C1FDFFFC",x"02200000",x"C1FDFFFC",x"02600006",x"40200000",x"C45C0000",x"C43C0004",x"C17DFFFC",x"00260000",x"03DC0010",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0010",x"C05C0004",x"C8240000",x"8A203D78",x"C07C0000",x"C0860018",x"C8240000",x"8E203D14",x"02A00000",x"82003D18",x"02A00001",x"82803D30",x"8E203D28",x"02800001",x"82003D2C",x"02800000",x"82003D34",x"008A0000",x"C0A60010",x"C82A0000",x"82803D44",x"82003D48",x"44202000",x"CC220000",x"C8240000",x"C43C0008",x"C17DFFFC",x"03DC0014",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0014",x"C03C0008",x"CC220004",x"82003D7C",x"CC020004",x"C05C0004",x"C8240004",x"8A203E04",x"C07C0000",x"C0860018",x"C8240004",x"8E203DA0",x"02A00000",x"82003DA4",x"02A00001",x"82803DBC",x"8E203DB4",x"02800001",x"82003DB8",x"02800000",x"82003DC0",x"008A0000",x"C0A60010",x"C82A0004",x"82803DD0",x"82003DD4",x"44202000",x"CC220008",x"C8240004",x"C43C0008",x"C17DFFFC",x"03DC0014",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0014",x"C03C0008",x"CC22000C",x"82003E08",x"CC02000C",x"C05C0004",x"C8240008",x"8A203E90",x"C07C0000",x"C0860018",x"C8240008",x"8E203E2C",x"02A00000",x"82003E30",x"02A00001",x"82803E48",x"8E203E40",x"02800001",x"82003E44",x"02800000",x"82003E4C",x"008A0000",x"C0660010",x"C8260008",x"82803E5C",x"82003E60",x"44202000",x"CC220010",x"C8240008",x"C43C0008",x"C17DFFFC",x"03DC0014",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0014",x"C03C0008",x"CC220014",x"82003E94",x"CC020014",x"C1FDFFFC",x"02600004",x"40200000",x"C45C0000",x"C43C0004",x"C17DFFFC",x"00260000",x"03DC0010",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0010",x"C05C0004",x"C8240000",x"C07C0000",x"C0860010",x"C8480000",x"48224000",x"C8440004",x"C0860010",x"C8680004",x"48446000",x"40224000",x"C8440008",x"C0460010",x"C8640008",x"48446000",x"40224000",x"8E023F10",x"CC020000",x"82004008",x"CC3C0008",x"C43C0010",x"C17DFFFC",x"03DC001C",x"037E000C",x"C57DFFFC",x"82000844",x"07DC001C",x"44202000",x"C03C0010",x"CC220000",x"C05C0000",x"C0640010",x"C8260000",x"C85C0008",x"CC3C0018",x"C17DFFFC",x"40204000",x"03DC0028",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0028",x"C85C0018",x"48242000",x"44202000",x"C03C0010",x"CC220004",x"C05C0000",x"C0640010",x"C8260004",x"C85C0008",x"CC3C0020",x"C17DFFFC",x"40204000",x"03DC0030",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0030",x"C85C0020",x"48242000",x"44202000",x"C03C0010",x"CC220008",x"C05C0000",x"C0440010",x"C8240008",x"C85C0008",x"CC3C0028",x"C17DFFFC",x"40204000",x"03DC0038",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0038",x"C85C0028",x"48242000",x"44202000",x"C03C0010",x"CC22000C",x"C1FDFFFC",x"02600005",x"40200000",x"C45C0000",x"C43C0004",x"C17DFFFC",x"00260000",x"03DC0010",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0010",x"C05C0004",x"C8240000",x"C8440004",x"C8640008",x"48822000",x"C07C0000",x"C0860010",x"C8A80000",x"4888A000",x"48A44000",x"C0860010",x"C8C80004",x"48AAC000",x"4088A000",x"48A66000",x"C0860010",x"C8C80008",x"48AAC000",x"4088A000",x"C086000C",x"828040CC",x"48A46000",x"C0860024",x"C8C80000",x"48AAC000",x"4088A000",x"48662000",x"C0860024",x"C8A80004",x"4866A000",x"40686000",x"48224000",x"C0860024",x"C8480008",x"48224000",x"40262000",x"820040D0",x"40208000",x"C8440000",x"C0860010",x"C8680000",x"48446000",x"44404000",x"C8640004",x"C0860010",x"C8880004",x"48668000",x"44606000",x"C8840008",x"C0860010",x"C8A80008",x"4888A000",x"44808000",x"CC220000",x"C086000C",x"CC3C0008",x"82804264",x"C8A40008",x"C0860024",x"C8C80004",x"48AAC000",x"C8C40004",x"C0860024",x"C8E80008",x"48CCE000",x"40AAC000",x"C8C00080",x"CC9C0010",x"CC7C0018",x"CCDC0020",x"C43C0028",x"CC5C0030",x"CCBC0038",x"C17DFFFC",x"4020C000",x"03DC0048",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0048",x"C85C0038",x"48242000",x"C85C0030",x"44242000",x"C03C0028",x"CC220004",x"C05C0004",x"C8240008",x"C07C0000",x"C0860024",x"C8480000",x"48224000",x"C8440000",x"C0860024",x"C8680008",x"48446000",x"40224000",x"C85C0020",x"CC3C0040",x"C17DFFFC",x"40204000",x"03DC0050",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0050",x"C85C0040",x"48242000",x"C85C0018",x"44242000",x"C03C0028",x"CC220008",x"C05C0004",x"C8240004",x"C07C0000",x"C0860024",x"C8480000",x"48224000",x"C8440000",x"C0460024",x"C8640004",x"48446000",x"40224000",x"C85C0020",x"CC3C0048",x"C17DFFFC",x"40204000",x"03DC0058",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0058",x"C85C0048",x"48242000",x"C85C0010",x"44242000",x"C03C0028",x"CC22000C",x"82004270",x"CC420004",x"CC620008",x"CC82000C",x"C83C0008",x"8A2042A0",x"C43C0028",x"C17DFFFC",x"03DC0058",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0058",x"C03C0028",x"CC220010",x"820042A0",x"C1FDFFFC",x"86404628",x"026000C8",x"22840220",x"D0868000",x"C0A20004",x"C0C20000",x"C0E80004",x"03000001",x"C43C0000",x"C47C0004",x"82F04350",x"03000002",x"82F04314",x"C4BC0008",x"C45C000C",x"C17DFFFC",x"00480000",x"002C0000",x"03DC0018",x"037E000C",x"C57DFFFC",x"8200400C",x"07DC0018",x"C05C000C",x"22640220",x"C09C0008",x"D4286000",x"8200434C",x"C4BC0008",x"C45C000C",x"C17DFFFC",x"00480000",x"002C0000",x"03DC0018",x"037E000C",x"C57DFFFC",x"82003E98",x"07DC0018",x"C05C000C",x"22640220",x"C09C0008",x"D4286000",x"82004388",x"C4BC0008",x"C45C000C",x"C17DFFFC",x"00480000",x"002C0000",x"03DC0018",x"037E000C",x"C57DFFFC",x"82003CC4",x"07DC0018",x"C05C000C",x"22640220",x"C09C0008",x"D4286000",x"06240001",x"86204624",x"22420220",x"C07C0004",x"D0464000",x"C09C0000",x"C0A80004",x"C0C80000",x"C0E40004",x"03000001",x"82F0442C",x"03000002",x"82F043F4",x"C4BC0010",x"C43C0014",x"C17DFFFC",x"002C0000",x"03DC0020",x"037E000C",x"C57DFFFC",x"8200400C",x"07DC0020",x"C05C0014",x"22640220",x"C09C0010",x"D4286000",x"82004428",x"C4BC0010",x"C43C0014",x"C17DFFFC",x"002C0000",x"03DC0020",x"037E000C",x"C57DFFFC",x"82003E98",x"07DC0020",x"C05C0014",x"22640220",x"C09C0010",x"D4286000",x"82004460",x"C4BC0010",x"C43C0014",x"C17DFFFC",x"002C0000",x"03DC0020",x"037E000C",x"C57DFFFC",x"82003CC4",x"07DC0020",x"C05C0014",x"22640220",x"C09C0010",x"D4286000",x"06240001",x"86204620",x"22420220",x"C07C0004",x"D0464000",x"C09C0000",x"C0A80004",x"C0C80000",x"C0E40004",x"03000001",x"82F04504",x"03000002",x"82F044CC",x"C4BC0018",x"C43C001C",x"C17DFFFC",x"002C0000",x"03DC0028",x"037E000C",x"C57DFFFC",x"8200400C",x"07DC0028",x"C05C001C",x"22640220",x"C09C0018",x"D4286000",x"82004500",x"C4BC0018",x"C43C001C",x"C17DFFFC",x"002C0000",x"03DC0028",x"037E000C",x"C57DFFFC",x"82003E98",x"07DC0028",x"C05C001C",x"22640220",x"C09C0018",x"D4286000",x"82004538",x"C4BC0018",x"C43C001C",x"C17DFFFC",x"002C0000",x"03DC0028",x"037E000C",x"C57DFFFC",x"82003CC4",x"07DC0028",x"C05C001C",x"22640220",x"C09C0018",x"D4286000",x"06240001",x"8620461C",x"22420220",x"C07C0004",x"D0464000",x"C07C0000",x"C0860004",x"C0A60000",x"C0C40004",x"02E00001",x"82CE45DC",x"02E00002",x"82CE45A4",x"C49C0020",x"C43C0024",x"C17DFFFC",x"002A0000",x"03DC0030",x"037E000C",x"C57DFFFC",x"8200400C",x"07DC0030",x"C05C0024",x"22640220",x"C09C0020",x"D4286000",x"820045D8",x"C49C0020",x"C43C0024",x"C17DFFFC",x"002A0000",x"03DC0030",x"037E000C",x"C57DFFFC",x"82003E98",x"07DC0030",x"C05C0024",x"22640220",x"C09C0020",x"D4286000",x"82004610",x"C49C0020",x"C43C0024",x"C17DFFFC",x"002A0000",x"03DC0030",x"037E000C",x"C57DFFFC",x"82003CC4",x"07DC0030",x"C05C0024",x"22640220",x"C09C0020",x"D4286000",x"06440001",x"C03C0000",x"820042A4",x"C1FDFFFC",x"C1FDFFFC",x"C1FDFFFC",x"C1FDFFFC",x"8640477C",x"026000C8",x"22840220",x"D0668000",x"C0860028",x"C0A60004",x"C8220000",x"C0C60014",x"C84C0000",x"44224000",x"CC280000",x"C8220004",x"C0C60014",x"C84C0004",x"44224000",x"CC280004",x"C8220008",x"C0C60014",x"C84C0008",x"44224000",x"CC280008",x"02C00002",x"82AC4740",x"02C00002",x"86CA4694",x"8200473C",x"C8280000",x"C8480004",x"C8680008",x"48822000",x"C0C60010",x"C8AC0000",x"4888A000",x"48A44000",x"C0C60010",x"C8CC0004",x"48AAC000",x"4088A000",x"48A66000",x"C0C60010",x"C8CC0008",x"48AAC000",x"4088A000",x"C0C6000C",x"82C04720",x"48A46000",x"C0C60024",x"C8CC0000",x"48AAC000",x"4088A000",x"48662000",x"C0C60024",x"C8AC0004",x"4866A000",x"40686000",x"48224000",x"C0660024",x"C8460008",x"48224000",x"40262000",x"82004724",x"40208000",x"02600003",x"82A64730",x"82004738",x"C84000A8",x"44224000",x"CC28000C",x"82004774",x"C0660010",x"C8280000",x"C8480004",x"C8680008",x"C8860000",x"48282000",x"C8860004",x"48484000",x"40224000",x"C8460008",x"48446000",x"40224000",x"CC28000C",x"06440001",x"8200462C",x"C1FDFFFC",x"48822000",x"C0420010",x"C8A40000",x"4888A000",x"48A44000",x"C0420010",x"C8C40004",x"48AAC000",x"4088A000",x"48A66000",x"C0420010",x"C8C40008",x"48AAC000",x"4088A000",x"C042000C",x"82404800",x"48A46000",x"C0420024",x"C8C40000",x"48AAC000",x"4088A000",x"48662000",x"C0420024",x"C8A40004",x"4866A000",x"40686000",x"48224000",x"C0420024",x"C8440008",x"48224000",x"40262000",x"82004804",x"40208000",x"C0420004",x"02600003",x"82464814",x"8200481C",x"C84000A8",x"44224000",x"C0220018",x"8E20482C",x"02400000",x"82004830",x"02400001",x"82204848",x"8E204840",x"02200001",x"82004844",x"02200000",x"8200484C",x"00240000",x"82204858",x"02200000",x"C1FDFFFC",x"02200001",x"C1FDFFFC",x"C0420014",x"C8840000",x"44228000",x"C0420014",x"C8840004",x"44448000",x"C0420014",x"C8840008",x"44668000",x"C0420004",x"02600001",x"8246497C",x"02600002",x"82464914",x"C43C0000",x"C17DFFFC",x"03DC000C",x"037E000C",x"C57DFFFC",x"82003344",x"07DC000C",x"C03C0000",x"C0420004",x"02600003",x"824648C8",x"820048D0",x"C84000A8",x"44224000",x"C0220018",x"8E2048E0",x"02400000",x"820048E4",x"02400001",x"822048FC",x"8E2048F4",x"02200001",x"820048F8",x"02200000",x"82004900",x"00240000",x"8220490C",x"02200000",x"C1FDFFFC",x"02200001",x"C1FDFFFC",x"C0420010",x"C8840000",x"48282000",x"C8840004",x"48484000",x"40224000",x"C8440008",x"48446000",x"40224000",x"C0220018",x"8E204948",x"02400000",x"8200494C",x"02400001",x"82204964",x"8E20495C",x"02200001",x"82004960",x"02200000",x"82004968",x"00240000",x"82204974",x"02200000",x"C1FDFFFC",x"02200001",x"C1FDFFFC",x"8E204984",x"82004988",x"44202000",x"C0420010",x"C8840000",x"8E28499C",x"02400000",x"820049E8",x"8E4049A8",x"40204000",x"820049AC",x"44204000",x"C0420010",x"C8440004",x"8E2449C0",x"02400000",x"820049E8",x"8E6049CC",x"40206000",x"820049D0",x"44206000",x"C0420010",x"C8440008",x"8E2449E4",x"02400000",x"820049E8",x"02400001",x"824049F4",x"C0220018",x"C1FDFFFC",x"C0220018",x"82204A04",x"02200000",x"C1FDFFFC",x"02200001",x"C1FDFFFC",x"22620220",x"D0646000",x"0280FFFF",x"82684E38",x"028000C8",x"22660220",x"D0686000",x"C0A60014",x"C88A0000",x"44828000",x"C0A60014",x"C8AA0004",x"44A4A000",x"C0A60014",x"C8CA0008",x"44C6C000",x"C0A60004",x"02C00001",x"CC7C0000",x"CC5C0008",x"CC3C0010",x"C49C0018",x"C45C001C",x"C43C0020",x"82AC4B0C",x"02C00002",x"82AC4AA4",x"C17DFFFC",x"00260000",x"4060C000",x"4040A000",x"40208000",x"03DC002C",x"037E000C",x"C57DFFFC",x"82004780",x"07DC002C",x"82004B08",x"C0A60010",x"C8EA0000",x"488E8000",x"C8EA0004",x"48AEA000",x"4088A000",x"C8AA0008",x"48AAC000",x"4088A000",x"C0660018",x"8E804AD8",x"02A00000",x"82004ADC",x"02A00001",x"82604AF4",x"8E804AEC",x"02600001",x"82004AF0",x"02600000",x"82004AF8",x"006A0000",x"82604B04",x"02200000",x"82004B08",x"02200001",x"82004B9C",x"8E804B14",x"82004B18",x"44808000",x"C0A60010",x"C8EA0000",x"8E8E4B2C",x"02A00000",x"82004B78",x"8EA04B38",x"4080A000",x"82004B3C",x"4480A000",x"C0A60010",x"C8AA0004",x"8E8A4B50",x"02A00000",x"82004B78",x"8EC04B5C",x"4080C000",x"82004B60",x"4480C000",x"C0A60010",x"C8AA0008",x"8E8A4B74",x"02A00000",x"82004B78",x"02A00001",x"82A04B88",x"C0660018",x"00260000",x"82004B9C",x"C0660018",x"82604B98",x"02200000",x"82004B9C",x"02200001",x"82204BA8",x"02200000",x"C1FDFFFC",x"C03C0020",x"02220001",x"22420220",x"C07C001C",x"D0464000",x"0280FFFF",x"82484E30",x"22440220",x"C09C0018",x"D0484000",x"C83C0010",x"C85C0008",x"C87C0000",x"C43C0024",x"C17DFFFC",x"00240000",x"03DC0030",x"037E000C",x"C57DFFFC",x"82004860",x"07DC0030",x"82204C08",x"02200000",x"C1FDFFFC",x"C03C0024",x"02220001",x"22420220",x"C07C001C",x"D0464000",x"0280FFFF",x"82484E28",x"22440220",x"C09C0018",x"D0484000",x"C0A40014",x"C82A0000",x"C85C0010",x"44242000",x"C0A40014",x"C86A0004",x"C89C0008",x"44686000",x"C0A40014",x"C8AA0008",x"C8DC0000",x"44ACA000",x"C0A40004",x"02C00001",x"C43C0028",x"82AC4D08",x"02C00002",x"82AC4CA0",x"C17DFFFC",x"00240000",x"40406000",x"4060A000",x"03DC0034",x"037E000C",x"C57DFFFC",x"82004780",x"07DC0034",x"82004D04",x"C0A40010",x"C8EA0000",x"482E2000",x"C8EA0004",x"486E6000",x"40226000",x"C86A0008",x"4866A000",x"40226000",x"C0440018",x"8E204CD4",x"02A00000",x"82004CD8",x"02A00001",x"82404CF0",x"8E204CE8",x"02400001",x"82004CEC",x"02400000",x"82004CF4",x"004A0000",x"82404D00",x"02200000",x"82004D04",x"02200001",x"82004D98",x"8E204D10",x"82004D14",x"44202000",x"C0A40010",x"C8EA0000",x"8E2E4D28",x"02A00000",x"82004D74",x"8E604D34",x"40206000",x"82004D38",x"44206000",x"C0A40010",x"C86A0004",x"8E264D4C",x"02A00000",x"82004D74",x"8EA04D58",x"4020A000",x"82004D5C",x"4420A000",x"C0A40010",x"C86A0008",x"8E264D70",x"02A00000",x"82004D74",x"02A00001",x"82A04D84",x"C0440018",x"00240000",x"82004D98",x"C0440018",x"82404D94",x"02200000",x"82004D98",x"02200001",x"82204DA4",x"02200000",x"C1FDFFFC",x"C03C0028",x"02220001",x"22420220",x"C07C001C",x"D0464000",x"0280FFFF",x"82484E20",x"22440220",x"C09C0018",x"D0484000",x"C83C0010",x"C85C0008",x"C87C0000",x"C43C002C",x"C17DFFFC",x"00240000",x"03DC0038",x"037E000C",x"C57DFFFC",x"82004860",x"07DC0038",x"82204E04",x"02200000",x"C1FDFFFC",x"C03C002C",x"02220001",x"C83C0010",x"C85C0008",x"C87C0000",x"C05C001C",x"82004A0C",x"02200001",x"C1FDFFFC",x"02200001",x"C1FDFFFC",x"02200001",x"C1FDFFFC",x"02200001",x"C1FDFFFC",x"22620220",x"D0646000",x"0280FFFF",x"8268527C",x"02800368",x"02A002B8",x"02C000C8",x"22E60220",x"D0ECE000",x"C82A0000",x"C10E0014",x"C8500000",x"44224000",x"C84A0004",x"C10E0014",x"C8700004",x"44446000",x"C86A0008",x"C10E0014",x"C8900008",x"44668000",x"C1080004",x"23260220",x"D1112000",x"C12E0004",x"03400001",x"C4BC0000",x"C45C0004",x"C43C0008",x"C4DC000C",x"C47C0010",x"83344F2C",x"02800002",x"83284EEC",x"C17DFFFC",x"00500000",x"002E0000",x"03DC001C",x"037E000C",x"C57DFFFC",x"82003A54",x"07DC001C",x"82004F28",x"C8900000",x"8E804EFC",x"02200000",x"82004F28",x"028002AC",x"C8900004",x"48282000",x"C8900008",x"48484000",x"40224000",x"C850000C",x"48446000",x"40224000",x"CC280000",x"02200001",x"82004F54",x"C0880000",x"C17DFFFC",x"00700000",x"00480000",x"002E0000",x"03DC001C",x"037E000C",x"C57DFFFC",x"8200389C",x"07DC001C",x"024002AC",x"C8240000",x"82204F78",x"C8400078",x"8E244F70",x"02200000",x"82004F74",x"02200001",x"82004F7C",x"02200000",x"8220524C",x"C8400074",x"40224000",x"022001D0",x"C8420000",x"48442000",x"C05C0000",x"C8640000",x"40446000",x"C8620004",x"48662000",x"C8840004",x"40668000",x"C8820008",x"48282000",x"C8840008",x"40228000",x"C05C0004",x"C0240000",x"0260FFFF",x"8226522C",x"22220220",x"C07C000C",x"D0262000",x"CC3C0018",x"CC7C0020",x"CC5C0028",x"C17DFFFC",x"41E06000",x"40602000",x"40204000",x"4041E000",x"03DC0038",x"037E000C",x"C57DFFFC",x"82004860",x"07DC0038",x"8220501C",x"02200000",x"82005228",x"C05C0004",x"C0240004",x"0260FFFF",x"82265224",x"22220220",x"C07C000C",x"D0262000",x"C0820014",x"C8280000",x"C85C0028",x"44242000",x"C0820014",x"C8680004",x"C89C0020",x"44686000",x"C0820014",x"C8A80008",x"C8DC0018",x"44ACA000",x"C0820004",x"02A00001",x"828A5108",x"02A00002",x"828A50A0",x"C17DFFFC",x"40406000",x"4060A000",x"03DC0038",x"037E000C",x"C57DFFFC",x"82004780",x"07DC0038",x"82005104",x"C0820010",x"C8E80000",x"482E2000",x"C8E80004",x"486E6000",x"40226000",x"C8680008",x"4866A000",x"40226000",x"C0220018",x"8E2050D4",x"02800000",x"820050D8",x"02800001",x"822050F0",x"8E2050E8",x"02200001",x"820050EC",x"02200000",x"820050F4",x"00280000",x"82205100",x"02200000",x"82005104",x"02200001",x"82005194",x"8E205110",x"82005114",x"44202000",x"C0820010",x"C8E80000",x"8E2E5128",x"02800000",x"82005174",x"8E605134",x"40206000",x"82005138",x"44206000",x"C0820010",x"C8680004",x"8E26514C",x"02800000",x"82005174",x"8EA05158",x"4020A000",x"8200515C",x"4420A000",x"C0820010",x"C8680008",x"8E265170",x"02800000",x"82005174",x"02800001",x"82805180",x"C0220018",x"82005194",x"C0220018",x"82205190",x"02200000",x"82005194",x"02200001",x"822051A0",x"02200000",x"82005220",x"C05C0004",x"C0240008",x"0260FFFF",x"8226521C",x"22220220",x"C07C000C",x"D0262000",x"C83C0028",x"C85C0020",x"C87C0018",x"C17DFFFC",x"03DC0038",x"037E000C",x"C57DFFFC",x"82004860",x"07DC0038",x"822051EC",x"02200000",x"82005218",x"02200003",x"C83C0028",x"C85C0020",x"C87C0018",x"C05C0004",x"C17DFFFC",x"03DC0038",x"037E000C",x"C57DFFFC",x"82004A0C",x"07DC0038",x"82005220",x"02200001",x"82005228",x"02200001",x"82005230",x"02200001",x"8220523C",x"02200001",x"C1FDFFFC",x"C03C0008",x"02220001",x"C05C0004",x"82004E40",x"C03C0010",x"22220220",x"C05C000C",x"D0242000",x"C0220018",x"82205274",x"C03C0008",x"02220001",x"C05C0004",x"82004E40",x"02200000",x"C1FDFFFC",x"02200000",x"C1FDFFFC",x"22620220",x"D0646000",x"0280FFFF",x"8268540C",x"028001E0",x"22660220",x"D0686000",x"02A00000",x"C49C0000",x"C45C0004",x"C43C0008",x"C17DFFFC",x"00460000",x"002A0000",x"03DC0014",x"037E000C",x"C57DFFFC",x"82004E40",x"07DC0014",x"822052DC",x"02200001",x"C1FDFFFC",x"C03C0008",x"02220001",x"22420220",x"C07C0004",x"D0464000",x"0280FFFF",x"82485404",x"22440220",x"C09C0000",x"D0484000",x"02A00000",x"C43C000C",x"C17DFFFC",x"002A0000",x"03DC0018",x"037E000C",x"C57DFFFC",x"82004E40",x"07DC0018",x"82205334",x"02200001",x"C1FDFFFC",x"C03C000C",x"02220001",x"22420220",x"C07C0004",x"D0464000",x"0280FFFF",x"824853FC",x"22440220",x"C09C0000",x"D0484000",x"02A00000",x"C43C0010",x"C17DFFFC",x"002A0000",x"03DC001C",x"037E000C",x"C57DFFFC",x"82004E40",x"07DC001C",x"8220538C",x"02200001",x"C1FDFFFC",x"C03C0010",x"02220001",x"22420220",x"C07C0004",x"D0464000",x"0280FFFF",x"824853F4",x"22440220",x"C09C0000",x"D0484000",x"02800000",x"C43C0014",x"C17DFFFC",x"00280000",x"03DC0020",x"037E000C",x"C57DFFFC",x"82004E40",x"07DC0020",x"822053E4",x"02200001",x"C1FDFFFC",x"C03C0014",x"02220001",x"C05C0004",x"82005284",x"02200000",x"C1FDFFFC",x"02200000",x"C1FDFFFC",x"02200000",x"C1FDFFFC",x"02200000",x"C1FDFFFC",x"22620220",x"D0646000",x"C0860000",x"02A0FFFF",x"828A57C0",x"02A00063",x"C47C0000",x"C45C0004",x"C43C0008",x"828A5678",x"02A00368",x"02C002B8",x"02E000C8",x"23080220",x"D0EF0000",x"C82C0000",x"C10E0014",x"C8500000",x"44224000",x"C84C0004",x"C10E0014",x"C8700004",x"44446000",x"C86C0008",x"C0CE0014",x"C88C0008",x"44668000",x"C0CA0004",x"22880220",x"D08C8000",x"C0CE0004",x"03000001",x"82D05504",x"02A00002",x"82CA54C4",x"C17DFFFC",x"00480000",x"002E0000",x"03DC0014",x"037E000C",x"C57DFFFC",x"82003A54",x"07DC0014",x"82005500",x"C8880000",x"8E8054D4",x"02200000",x"82005500",x"02A002AC",x"C8880004",x"48282000",x"C8880008",x"48484000",x"40224000",x"C848000C",x"48446000",x"40224000",x"CC2A0000",x"02200001",x"8200552C",x"C0AA0000",x"C17DFFFC",x"00680000",x"004A0000",x"002E0000",x"03DC0014",x"037E000C",x"C57DFFFC",x"8200389C",x"07DC0014",x"82205670",x"022002AC",x"C8220000",x"C8400070",x"8E245548",x"02200000",x"8200566C",x"C03C0000",x"C0420004",x"0260FFFF",x"82465658",x"026001E0",x"22440220",x"D0464000",x"02800000",x"C47C000C",x"C17DFFFC",x"00280000",x"03DC0018",x"037E000C",x"C57DFFFC",x"82004E40",x"07DC0018",x"82205594",x"02200001",x"82005654",x"C03C0000",x"C0420008",x"0260FFFF",x"82465650",x"22440220",x"C07C000C",x"D0464000",x"02800000",x"C17DFFFC",x"00280000",x"03DC0018",x"037E000C",x"C57DFFFC",x"82004E40",x"07DC0018",x"822055DC",x"02200001",x"8200564C",x"C03C0000",x"C042000C",x"0260FFFF",x"82465648",x"22440220",x"C07C000C",x"D0464000",x"02600000",x"C17DFFFC",x"00260000",x"03DC0018",x"037E000C",x"C57DFFFC",x"82004E40",x"07DC0018",x"82205624",x"02200001",x"82005644",x"02200004",x"C05C0000",x"C17DFFFC",x"03DC0018",x"037E000C",x"C57DFFFC",x"82005284",x"07DC0018",x"8200564C",x"02200000",x"82005654",x"02200000",x"8200565C",x"02200000",x"82205668",x"02200001",x"8200566C",x"02200000",x"82005674",x"02200000",x"8200567C",x"02200001",x"822057B0",x"C03C0000",x"C0420004",x"0260FFFF",x"82465790",x"026001E0",x"22440220",x"D0464000",x"02800000",x"C47C0010",x"C17DFFFC",x"00280000",x"03DC001C",x"037E000C",x"C57DFFFC",x"82004E40",x"07DC001C",x"822056CC",x"02200001",x"8200578C",x"C03C0000",x"C0420008",x"0260FFFF",x"82465788",x"22440220",x"C07C0010",x"D0464000",x"02800000",x"C17DFFFC",x"00280000",x"03DC001C",x"037E000C",x"C57DFFFC",x"82004E40",x"07DC001C",x"82205714",x"02200001",x"82005784",x"C03C0000",x"C042000C",x"0260FFFF",x"82465780",x"22440220",x"C07C0010",x"D0464000",x"02600000",x"C17DFFFC",x"00260000",x"03DC001C",x"037E000C",x"C57DFFFC",x"82004E40",x"07DC001C",x"8220575C",x"02200001",x"8200577C",x"02200004",x"C05C0000",x"C17DFFFC",x"03DC001C",x"037E000C",x"C57DFFFC",x"82005284",x"07DC001C",x"82005784",x"02200000",x"8200578C",x"02200000",x"82005794",x"02200000",x"822057A0",x"02200001",x"C1FDFFFC",x"C03C0008",x"02220001",x"C05C0004",x"82005414",x"C03C0008",x"02220001",x"C05C0004",x"82005414",x"02200000",x"C1FDFFFC",x"22820220",x"D0848000",x"02A0FFFF",x"828A5CD8",x"02A0030C",x"02C000C8",x"22E80220",x"D0ECE000",x"C82A0000",x"C10E0014",x"C8500000",x"44224000",x"C84A0004",x"C10E0014",x"C8700004",x"44446000",x"C86A0008",x"C10E0014",x"C8900008",x"44668000",x"C10E0004",x"03200001",x"C4BC0000",x"C47C0004",x"C45C0008",x"C43C000C",x"C4DC0010",x"C49C0014",x"8312588C",x"03200002",x"83125868",x"C17DFFFC",x"00460000",x"002E0000",x"03DC0020",x"037E000C",x"C57DFFFC",x"820034A0",x"07DC0020",x"82005888",x"C17DFFFC",x"00460000",x"002E0000",x"03DC0020",x"037E000C",x"C57DFFFC",x"820032A4",x"07DC0020",x"8200596C",x"03000000",x"03200001",x"03400002",x"CC3C0018",x"CC7C0020",x"CC5C0028",x"C4FC0030",x"C17DFFFC",x"00B40000",x"00920000",x"00460000",x"002E0000",x"00700000",x"03DC003C",x"037E000C",x"C57DFFFC",x"8200317C",x"07DC003C",x"822058E0",x"02200001",x"8200596C",x"02600001",x"02800002",x"02A00000",x"C83C0028",x"C85C0020",x"C87C0018",x"C03C0030",x"C05C0004",x"C17DFFFC",x"03DC003C",x"037E000C",x"C57DFFFC",x"8200317C",x"07DC003C",x"82205924",x"02200002",x"8200596C",x"02600002",x"02800000",x"02A00001",x"C83C0020",x"C85C0018",x"C87C0028",x"C03C0030",x"C05C0004",x"C17DFFFC",x"03DC003C",x"037E000C",x"C57DFFFC",x"8200317C",x"07DC003C",x"82205968",x"02200003",x"8200596C",x"02200000",x"82205CA8",x"024002AC",x"C8240000",x"8E025980",x"82005C94",x"024002B4",x"C8440000",x"8E245990",x"82005C94",x"C8400074",x"40224000",x"C07C0004",x"C8460000",x"48442000",x"C09C0000",x"C8680000",x"40446000",x"C8660004",x"48662000",x"C8880004",x"40668000",x"C8860008",x"48882000",x"C8A80008",x"4088A000",x"C09C0008",x"C0A80000",x"02C0FFFF",x"C43C0034",x"CC9C0038",x"CC7C0040",x"CC5C0048",x"C45C0050",x"CC3C0058",x"82AC5C48",x"22AA0220",x"C0DC0010",x"D0ACA000",x"C17DFFFC",x"002A0000",x"40204000",x"40406000",x"40608000",x"03DC0068",x"037E000C",x"C57DFFFC",x"82004860",x"07DC0068",x"82205A38",x"02200000",x"82005C44",x"C05C0008",x"C0240004",x"0260FFFF",x"82265C40",x"22220220",x"C07C0010",x"D0262000",x"C0820014",x"C8280000",x"C85C0048",x"44242000",x"C0820014",x"C8680004",x"C89C0040",x"44686000",x"C0820014",x"C8A80008",x"C8DC0038",x"44ACA000",x"C0820004",x"02A00001",x"828A5B24",x"02A00002",x"828A5ABC",x"C17DFFFC",x"40406000",x"4060A000",x"03DC0068",x"037E000C",x"C57DFFFC",x"82004780",x"07DC0068",x"82005B20",x"C0820010",x"C8E80000",x"482E2000",x"C8E80004",x"486E6000",x"40226000",x"C8680008",x"4866A000",x"40226000",x"C0220018",x"8E205AF0",x"02800000",x"82005AF4",x"02800001",x"82205B0C",x"8E205B04",x"02200001",x"82005B08",x"02200000",x"82005B10",x"00280000",x"82205B1C",x"02200000",x"82005B20",x"02200001",x"82005BB0",x"8E205B2C",x"82005B30",x"44202000",x"C0820010",x"C8E80000",x"8E2E5B44",x"02800000",x"82005B90",x"8E605B50",x"40206000",x"82005B54",x"44206000",x"C0820010",x"C8680004",x"8E265B68",x"02800000",x"82005B90",x"8EA05B74",x"4020A000",x"82005B78",x"4420A000",x"C0820010",x"C8680008",x"8E265B8C",x"02800000",x"82005B90",x"02800001",x"82805B9C",x"C0220018",x"82005BB0",x"C0220018",x"82205BAC",x"02200000",x"82005BB0",x"02200001",x"82205BBC",x"02200000",x"82005C3C",x"C05C0008",x"C0240008",x"0260FFFF",x"82265C38",x"22220220",x"C07C0010",x"D0262000",x"C83C0048",x"C85C0040",x"C87C0038",x"C17DFFFC",x"03DC0068",x"037E000C",x"C57DFFFC",x"82004860",x"07DC0068",x"82205C08",x"02200000",x"82005C34",x"02200003",x"C83C0048",x"C85C0040",x"C87C0038",x"C05C0008",x"C17DFFFC",x"03DC0068",x"037E000C",x"C57DFFFC",x"82004A0C",x"07DC0068",x"82005C3C",x"02200001",x"82005C44",x"02200001",x"82005C4C",x"02200001",x"82205C94",x"C03C0050",x"C83C0058",x"CC220000",x"022002B8",x"C83C0048",x"CC220000",x"C83C0040",x"CC220004",x"C83C0038",x"CC220008",x"022002C4",x"C05C0014",x"C4420000",x"022002B0",x"C05C0034",x"C4420000",x"82005C94",x"C03C000C",x"02220001",x"C05C0008",x"C07C0004",x"820057C8",x"C03C0014",x"22220220",x"C05C0010",x"D0242000",x"C0220018",x"82205CD4",x"C03C000C",x"02220001",x"C05C0008",x"C07C0004",x"820057C8",x"C1FDFFFC",x"C1FDFFFC",x"22820220",x"D0848000",x"02A0FFFF",x"828A5E48",x"02A001E0",x"22880220",x"D08A8000",x"02C00000",x"C47C0000",x"C4BC0004",x"C45C0008",x"C43C000C",x"C17DFFFC",x"00480000",x"002C0000",x"03DC0018",x"037E000C",x"C57DFFFC",x"820057C8",x"07DC0018",x"C03C000C",x"02220001",x"22420220",x"C07C0008",x"D0464000",x"0280FFFF",x"82485E44",x"22440220",x"C09C0004",x"D0484000",x"02A00000",x"C0DC0000",x"C43C0010",x"C17DFFFC",x"006C0000",x"002A0000",x"03DC001C",x"037E000C",x"C57DFFFC",x"820057C8",x"07DC001C",x"C03C0010",x"02220001",x"22420220",x"C07C0008",x"D0464000",x"0280FFFF",x"82485E40",x"22440220",x"C09C0004",x"D0484000",x"02A00000",x"C0DC0000",x"C43C0014",x"C17DFFFC",x"006C0000",x"002A0000",x"03DC0020",x"037E000C",x"C57DFFFC",x"820057C8",x"07DC0020",x"C03C0014",x"02220001",x"22420220",x"C07C0008",x"D0464000",x"0280FFFF",x"82485E3C",x"22440220",x"C09C0004",x"D0484000",x"02800000",x"C0BC0000",x"C43C0018",x"C17DFFFC",x"006A0000",x"00280000",x"03DC0024",x"037E000C",x"C57DFFFC",x"820057C8",x"07DC0024",x"C03C0018",x"02220001",x"C05C0008",x"C07C0000",x"82005CDC",x"C1FDFFFC",x"C1FDFFFC",x"C1FDFFFC",x"C1FDFFFC",x"22820220",x"D0848000",x"C0A80000",x"02C0FFFF",x"82AC6420",x"02C00063",x"C47C0000",x"C45C0004",x"C43C0008",x"82AC6118",x"02C0030C",x"02E000C8",x"22AA0220",x"D0AEA000",x"C82C0000",x"C0EA0014",x"C84E0000",x"44224000",x"C84C0004",x"C0EA0014",x"C86E0004",x"44446000",x"C86C0008",x"C0CA0014",x"C88C0008",x"44668000",x"C0CA0004",x"02E00001",x"C49C000C",x"82CE5F14",x"02E00002",x"82CE5EF0",x"C17DFFFC",x"00460000",x"002A0000",x"03DC0018",x"037E000C",x"C57DFFFC",x"820034A0",x"07DC0018",x"82005F10",x"C17DFFFC",x"00460000",x"002A0000",x"03DC0018",x"037E000C",x"C57DFFFC",x"820032A4",x"07DC0018",x"82005FF4",x"02C00000",x"02E00001",x"03000002",x"CC3C0010",x"CC7C0018",x"CC5C0020",x"C4BC0028",x"C17DFFFC",x"008E0000",x"00460000",x"002A0000",x"00B00000",x"006C0000",x"03DC0034",x"037E000C",x"C57DFFFC",x"8200317C",x"07DC0034",x"82205F68",x"02200001",x"82005FF4",x"02600001",x"02800002",x"02A00000",x"C83C0020",x"C85C0018",x"C87C0010",x"C03C0028",x"C05C0000",x"C17DFFFC",x"03DC0034",x"037E000C",x"C57DFFFC",x"8200317C",x"07DC0034",x"82205FAC",x"02200002",x"82005FF4",x"02600002",x"02800000",x"02A00001",x"C83C0018",x"C85C0010",x"C87C0020",x"C03C0028",x"C05C0000",x"C17DFFFC",x"03DC0034",x"037E000C",x"C57DFFFC",x"8200317C",x"07DC0034",x"82205FF0",x"02200003",x"82005FF4",x"02200000",x"82206114",x"022002AC",x"C8220000",x"022002B4",x"C8420000",x"8E246010",x"82006110",x"C03C000C",x"C0420004",x"0260FFFF",x"82466110",x"026001E0",x"22440220",x"D0464000",x"02800000",x"C0BC0000",x"C47C002C",x"C17DFFFC",x"006A0000",x"00280000",x"03DC0038",x"037E000C",x"C57DFFFC",x"820057C8",x"07DC0038",x"C03C000C",x"C0420008",x"0260FFFF",x"8246610C",x"22440220",x"C07C002C",x"D0464000",x"02800000",x"C0BC0000",x"C17DFFFC",x"006A0000",x"00280000",x"03DC0038",x"037E000C",x"C57DFFFC",x"820057C8",x"07DC0038",x"C03C000C",x"C042000C",x"0260FFFF",x"82466108",x"22440220",x"C07C002C",x"D0464000",x"02600000",x"C09C0000",x"C17DFFFC",x"00260000",x"00680000",x"03DC0038",x"037E000C",x"C57DFFFC",x"820057C8",x"07DC0038",x"02200004",x"C05C000C",x"C07C0000",x"C17DFFFC",x"03DC0038",x"037E000C",x"C57DFFFC",x"82005CDC",x"07DC0038",x"82006108",x"8200610C",x"82006110",x"82006114",x"82006214",x"C0A80004",x"02C0FFFF",x"82AC6214",x"02C001E0",x"22AA0220",x"D0ACA000",x"02E00000",x"C4DC0030",x"C49C000C",x"C17DFFFC",x"004A0000",x"002E0000",x"03DC003C",x"037E000C",x"C57DFFFC",x"820057C8",x"07DC003C",x"C03C000C",x"C0420008",x"0260FFFF",x"82466210",x"22440220",x"C07C0030",x"D0464000",x"02800000",x"C0BC0000",x"C17DFFFC",x"006A0000",x"00280000",x"03DC003C",x"037E000C",x"C57DFFFC",x"820057C8",x"07DC003C",x"C03C000C",x"C042000C",x"0260FFFF",x"8246620C",x"22440220",x"C07C0030",x"D0464000",x"02600000",x"C09C0000",x"C17DFFFC",x"00260000",x"00680000",x"03DC003C",x"037E000C",x"C57DFFFC",x"820057C8",x"07DC003C",x"02200004",x"C05C000C",x"C07C0000",x"C17DFFFC",x"03DC003C",x"037E000C",x"C57DFFFC",x"82005CDC",x"07DC003C",x"8200620C",x"82006210",x"82006214",x"C03C0008",x"02220001",x"22420220",x"C07C0004",x"D0464000",x"C0840000",x"02A0FFFF",x"828A641C",x"02A00063",x"C43C0034",x"828A634C",x"02A0030C",x"C0DC0000",x"C45C0038",x"C17DFFFC",x"006A0000",x"004C0000",x"00280000",x"03DC0044",x"037E000C",x"C57DFFFC",x"820036D4",x"07DC0044",x"82206348",x"022002AC",x"C8220000",x"022002B4",x"C8420000",x"8E24628C",x"82006344",x"C03C0038",x"C0420004",x"0260FFFF",x"82466344",x"026001E0",x"22440220",x"D0464000",x"02800000",x"C0BC0000",x"C47C003C",x"C17DFFFC",x"006A0000",x"00280000",x"03DC0048",x"037E000C",x"C57DFFFC",x"820057C8",x"07DC0048",x"C03C0038",x"C0420008",x"0260FFFF",x"82466340",x"22440220",x"C07C003C",x"D0464000",x"02600000",x"C09C0000",x"C17DFFFC",x"00260000",x"00680000",x"03DC0048",x"037E000C",x"C57DFFFC",x"820057C8",x"07DC0048",x"02200003",x"C05C0038",x"C07C0000",x"C17DFFFC",x"03DC0048",x"037E000C",x"C57DFFFC",x"82005CDC",x"07DC0048",x"82006340",x"82006344",x"82006348",x"82006408",x"C0840004",x"02A0FFFF",x"828A6408",x"02A001E0",x"22880220",x"D08A8000",x"02C00000",x"C0FC0000",x"C4BC0040",x"C45C0038",x"C17DFFFC",x"006E0000",x"00480000",x"002C0000",x"03DC004C",x"037E000C",x"C57DFFFC",x"820057C8",x"07DC004C",x"C03C0038",x"C0420008",x"0260FFFF",x"82466404",x"22440220",x"C07C0040",x"D0464000",x"02600000",x"C09C0000",x"C17DFFFC",x"00260000",x"00680000",x"03DC004C",x"037E000C",x"C57DFFFC",x"820057C8",x"07DC004C",x"02200003",x"C05C0038",x"C07C0000",x"C17DFFFC",x"03DC004C",x"037E000C",x"C57DFFFC",x"82005CDC",x"07DC004C",x"82006404",x"82006408",x"C03C0034",x"02220001",x"C05C0004",x"C07C0000",x"82005E4C",x"C1FDFFFC",x"C1FDFFFC",x"C0860000",x"22A20220",x"D0A4A000",x"02C0FFFF",x"82AC6874",x"02C000C8",x"22EA0220",x"D0ECE000",x"C10E0028",x"C8300000",x"C8500004",x"C8700008",x"C1260004",x"234A0220",x"D1334000",x"C14E0004",x"C49C0000",x"02800001",x"C47C0004",x"C45C0008",x"C43C000C",x"C4DC0010",x"C4BC0014",x"834864E0",x"02800002",x"834864B4",x"C17DFFFC",x"00700000",x"00520000",x"002E0000",x"03DC0020",x"037E000C",x"C57DFFFC",x"82003BD4",x"07DC0020",x"820064DC",x"C8320000",x"8E2064C4",x"02200000",x"820064DC",x"028002AC",x"C8320000",x"C850000C",x"48224000",x"CC280000",x"02200001",x"82006508",x"C0860000",x"C17DFFFC",x"00720000",x"00480000",x"002E0000",x"03DC0020",x"037E000C",x"C57DFFFC",x"8200389C",x"07DC0020",x"82206844",x"024002AC",x"C8240000",x"8E02651C",x"82006830",x"024002B4",x"C8440000",x"8E24652C",x"82006830",x"C8400074",x"40224000",x"C07C0000",x"C8460000",x"48442000",x"02800318",x"C8680000",x"40446000",x"C8660004",x"48662000",x"C8880004",x"40668000",x"C8860008",x"48882000",x"C8A80008",x"4088A000",x"C07C0008",x"C0860000",x"02A0FFFF",x"C43C0018",x"CC9C0020",x"CC7C0028",x"CC5C0030",x"C45C0038",x"CC3C0040",x"828A67E4",x"22880220",x"C0BC0010",x"D08A8000",x"C17DFFFC",x"00280000",x"40204000",x"40406000",x"40608000",x"03DC0050",x"037E000C",x"C57DFFFC",x"82004860",x"07DC0050",x"822065D4",x"02200000",x"820067E0",x"C05C0008",x"C0240004",x"0260FFFF",x"822667DC",x"22220220",x"C07C0010",x"D0262000",x"C0820014",x"C8280000",x"C85C0030",x"44242000",x"C0820014",x"C8680004",x"C89C0028",x"44686000",x"C0820014",x"C8A80008",x"C8DC0020",x"44ACA000",x"C0820004",x"02A00001",x"828A66C0",x"02A00002",x"828A6658",x"C17DFFFC",x"40406000",x"4060A000",x"03DC0050",x"037E000C",x"C57DFFFC",x"82004780",x"07DC0050",x"820066BC",x"C0820010",x"C8E80000",x"482E2000",x"C8E80004",x"486E6000",x"40226000",x"C8680008",x"4866A000",x"40226000",x"C0220018",x"8E20668C",x"02800000",x"82006690",x"02800001",x"822066A8",x"8E2066A0",x"02200001",x"820066A4",x"02200000",x"820066AC",x"00280000",x"822066B8",x"02200000",x"820066BC",x"02200001",x"8200674C",x"8E2066C8",x"820066CC",x"44202000",x"C0820010",x"C8E80000",x"8E2E66E0",x"02800000",x"8200672C",x"8E6066EC",x"40206000",x"820066F0",x"44206000",x"C0820010",x"C8680004",x"8E266704",x"02800000",x"8200672C",x"8EA06710",x"4020A000",x"82006714",x"4420A000",x"C0820010",x"C8680008",x"8E266728",x"02800000",x"8200672C",x"02800001",x"82806738",x"C0220018",x"8200674C",x"C0220018",x"82206748",x"02200000",x"8200674C",x"02200001",x"82206758",x"02200000",x"820067D8",x"C05C0008",x"C0240008",x"0260FFFF",x"822667D4",x"22220220",x"C07C0010",x"D0262000",x"C83C0030",x"C85C0028",x"C87C0020",x"C17DFFFC",x"03DC0050",x"037E000C",x"C57DFFFC",x"82004860",x"07DC0050",x"822067A4",x"02200000",x"820067D0",x"02200003",x"C83C0030",x"C85C0028",x"C87C0020",x"C05C0008",x"C17DFFFC",x"03DC0050",x"037E000C",x"C57DFFFC",x"82004A0C",x"07DC0050",x"820067D8",x"02200001",x"820067E0",x"02200001",x"820067E8",x"02200001",x"82206830",x"C03C0038",x"C83C0040",x"CC220000",x"022002B8",x"C83C0030",x"CC220000",x"C83C0028",x"CC220004",x"C83C0020",x"CC220008",x"022002C4",x"C05C0014",x"C4420000",x"022002B0",x"C05C0018",x"C4420000",x"82006830",x"C03C000C",x"02220001",x"C05C0008",x"C07C0004",x"82006424",x"C03C0014",x"22220220",x"C05C0010",x"D0242000",x"C0220018",x"82206870",x"C03C000C",x"02220001",x"C05C0008",x"C07C0004",x"82006424",x"C1FDFFFC",x"C1FDFFFC",x"22820220",x"D0848000",x"02A0FFFF",x"828A69E4",x"02A001E0",x"22880220",x"D08A8000",x"02C00000",x"C47C0000",x"C4BC0004",x"C45C0008",x"C43C000C",x"C17DFFFC",x"00480000",x"002C0000",x"03DC0018",x"037E000C",x"C57DFFFC",x"82006424",x"07DC0018",x"C03C000C",x"02220001",x"22420220",x"C07C0008",x"D0464000",x"0280FFFF",x"824869E0",x"22440220",x"C09C0004",x"D0484000",x"02A00000",x"C0DC0000",x"C43C0010",x"C17DFFFC",x"006C0000",x"002A0000",x"03DC001C",x"037E000C",x"C57DFFFC",x"82006424",x"07DC001C",x"C03C0010",x"02220001",x"22420220",x"C07C0008",x"D0464000",x"0280FFFF",x"824869DC",x"22440220",x"C09C0004",x"D0484000",x"02A00000",x"C0DC0000",x"C43C0014",x"C17DFFFC",x"006C0000",x"002A0000",x"03DC0020",x"037E000C",x"C57DFFFC",x"82006424",x"07DC0020",x"C03C0014",x"02220001",x"22420220",x"C07C0008",x"D0464000",x"0280FFFF",x"824869D8",x"22440220",x"C09C0004",x"D0484000",x"02800000",x"C0BC0000",x"C43C0018",x"C17DFFFC",x"006A0000",x"00280000",x"03DC0024",x"037E000C",x"C57DFFFC",x"82006424",x"07DC0024",x"C03C0018",x"02220001",x"C05C0008",x"C07C0000",x"82006878",x"C1FDFFFC",x"C1FDFFFC",x"C1FDFFFC",x"C1FDFFFC",x"22820220",x"D0848000",x"C0A80000",x"02C0FFFF",x"82AC6F88",x"02C00063",x"C47C0000",x"C45C0004",x"C43C0008",x"82AC6BF0",x"02C000C8",x"22EA0220",x"D0CCE000",x"C0EC0028",x"C82E0000",x"C84E0004",x"C86E0008",x"C1060004",x"22AA0220",x"D0B0A000",x"C10C0004",x"03200001",x"C49C000C",x"83126AA4",x"03200002",x"83126A78",x"C17DFFFC",x"006E0000",x"004A0000",x"002C0000",x"03DC0018",x"037E000C",x"C57DFFFC",x"82003BD4",x"07DC0018",x"82006AA0",x"C82A0000",x"8E206A88",x"02200000",x"82006AA0",x"02C002AC",x"C82A0000",x"C84E000C",x"48224000",x"CC2C0000",x"02200001",x"82006ACC",x"C0E60000",x"C17DFFFC",x"006A0000",x"004E0000",x"002C0000",x"03DC0018",x"037E000C",x"C57DFFFC",x"8200389C",x"07DC0018",x"82206BEC",x"022002AC",x"C8220000",x"022002B4",x"C8420000",x"8E246AE8",x"82006BE8",x"C03C000C",x"C0420004",x"0260FFFF",x"82466BE8",x"026001E0",x"22440220",x"D0464000",x"02800000",x"C0BC0000",x"C47C0010",x"C17DFFFC",x"006A0000",x"00280000",x"03DC001C",x"037E000C",x"C57DFFFC",x"82006424",x"07DC001C",x"C03C000C",x"C0420008",x"0260FFFF",x"82466BE4",x"22440220",x"C07C0010",x"D0464000",x"02800000",x"C0BC0000",x"C17DFFFC",x"006A0000",x"00280000",x"03DC001C",x"037E000C",x"C57DFFFC",x"82006424",x"07DC001C",x"C03C000C",x"C042000C",x"0260FFFF",x"82466BE0",x"22440220",x"C07C0010",x"D0464000",x"02600000",x"C09C0000",x"C17DFFFC",x"00260000",x"00680000",x"03DC001C",x"037E000C",x"C57DFFFC",x"82006424",x"07DC001C",x"02200004",x"C05C000C",x"C07C0000",x"C17DFFFC",x"03DC001C",x"037E000C",x"C57DFFFC",x"82006878",x"07DC001C",x"82006BE0",x"82006BE4",x"82006BE8",x"82006BEC",x"82006CEC",x"C0A80004",x"02C0FFFF",x"82AC6CEC",x"02C001E0",x"22AA0220",x"D0ACA000",x"02E00000",x"C4DC0014",x"C49C000C",x"C17DFFFC",x"004A0000",x"002E0000",x"03DC0020",x"037E000C",x"C57DFFFC",x"82006424",x"07DC0020",x"C03C000C",x"C0420008",x"0260FFFF",x"82466CE8",x"22440220",x"C07C0014",x"D0464000",x"02800000",x"C0BC0000",x"C17DFFFC",x"006A0000",x"00280000",x"03DC0020",x"037E000C",x"C57DFFFC",x"82006424",x"07DC0020",x"C03C000C",x"C042000C",x"0260FFFF",x"82466CE4",x"22440220",x"C07C0014",x"D0464000",x"02600000",x"C09C0000",x"C17DFFFC",x"00260000",x"00680000",x"03DC0020",x"037E000C",x"C57DFFFC",x"82006424",x"07DC0020",x"02200004",x"C05C000C",x"C07C0000",x"C17DFFFC",x"03DC0020",x"037E000C",x"C57DFFFC",x"82006878",x"07DC0020",x"82006CE4",x"82006CE8",x"82006CEC",x"C03C0008",x"02220001",x"22420220",x"C07C0004",x"D0464000",x"C0840000",x"02A0FFFF",x"828A6F84",x"02A00063",x"C43C0018",x"828A6EB4",x"02A000C8",x"22C80220",x"D0AAC000",x"C0CA0028",x"C82C0000",x"C84C0004",x"C86C0008",x"C0FC0000",x"C10E0004",x"22880220",x"D0908000",x"C10A0004",x"03200001",x"C45C001C",x"83126DB0",x"03200002",x"83126D84",x"C17DFFFC",x"006C0000",x"00480000",x"002A0000",x"03DC0028",x"037E000C",x"C57DFFFC",x"82003BD4",x"07DC0028",x"82006DAC",x"C8280000",x"8E206D94",x"02200000",x"82006DAC",x"02A002AC",x"C8280000",x"C84C000C",x"48224000",x"CC2A0000",x"02200001",x"82006DD8",x"C0CE0000",x"C17DFFFC",x"00680000",x"004C0000",x"002A0000",x"03DC0028",x"037E000C",x"C57DFFFC",x"8200389C",x"07DC0028",x"82206EB0",x"022002AC",x"C8220000",x"022002B4",x"C8420000",x"8E246DF4",x"82006EAC",x"C03C001C",x"C0420004",x"0260FFFF",x"82466EAC",x"026001E0",x"22440220",x"D0464000",x"02800000",x"C0BC0000",x"C47C0020",x"C17DFFFC",x"006A0000",x"00280000",x"03DC002C",x"037E000C",x"C57DFFFC",x"82006424",x"07DC002C",x"C03C001C",x"C0420008",x"0260FFFF",x"82466EA8",x"22440220",x"C07C0020",x"D0464000",x"02600000",x"C09C0000",x"C17DFFFC",x"00260000",x"00680000",x"03DC002C",x"037E000C",x"C57DFFFC",x"82006424",x"07DC002C",x"02200003",x"C05C001C",x"C07C0000",x"C17DFFFC",x"03DC002C",x"037E000C",x"C57DFFFC",x"82006878",x"07DC002C",x"82006EA8",x"82006EAC",x"82006EB0",x"82006F70",x"C0840004",x"02A0FFFF",x"828A6F70",x"02A001E0",x"22880220",x"D08A8000",x"02C00000",x"C0FC0000",x"C4BC0024",x"C45C001C",x"C17DFFFC",x"006E0000",x"00480000",x"002C0000",x"03DC0030",x"037E000C",x"C57DFFFC",x"82006424",x"07DC0030",x"C03C001C",x"C0420008",x"0260FFFF",x"82466F6C",x"22440220",x"C07C0024",x"D0464000",x"02600000",x"C09C0000",x"C17DFFFC",x"00260000",x"00680000",x"03DC0030",x"037E000C",x"C57DFFFC",x"82006424",x"07DC0030",x"02200003",x"C05C001C",x"C07C0000",x"C17DFFFC",x"03DC0030",x"037E000C",x"C57DFFFC",x"82006878",x"07DC0030",x"82006F6C",x"82006F70",x"C03C0018",x"02220001",x"C05C0004",x"C07C0000",x"820069E8",x"C1FDFFFC",x"C1FDFFFC",x"024002B8",x"C8240000",x"C0620014",x"C8460000",x"44224000",x"C8440004",x"C0620014",x"C8660004",x"44446000",x"C8640008",x"C0420014",x"C8840008",x"44668000",x"C0420010",x"C8840000",x"48828000",x"C0420010",x"C8A40004",x"48A4A000",x"C0420010",x"C8C40008",x"48C6C000",x"C042000C",x"C43C0000",x"82407138",x"024002C8",x"C0620024",x"C8E60008",x"48E4E000",x"C0620024",x"C9060004",x"49070000",x"40EF0000",x"C9000080",x"CCDC0008",x"CC5C0010",x"CCBC0018",x"CD1C0020",x"CC7C0028",x"CC3C0030",x"C45C0038",x"CC9C0040",x"CCFC0048",x"C17DFFFC",x"40210000",x"03DC0058",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0058",x"C85C0048",x"48242000",x"C85C0040",x"40242000",x"C03C0038",x"CC220000",x"C05C0000",x"C0640024",x"C8260008",x"C85C0030",x"48242000",x"C0640024",x"C8660000",x"C89C0028",x"48686000",x"40226000",x"C87C0020",x"CC3C0050",x"C17DFFFC",x"40206000",x"03DC0060",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0060",x"C85C0050",x"48242000",x"C85C0018",x"40242000",x"C03C0038",x"CC220004",x"C05C0000",x"C0640024",x"C8260004",x"C85C0030",x"48242000",x"C0640024",x"C8460000",x"C87C0010",x"48464000",x"40224000",x"C85C0020",x"CC3C0058",x"C17DFFFC",x"40204000",x"03DC0068",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0068",x"C85C0058",x"48242000",x"C85C0008",x"40242000",x"C03C0038",x"CC220008",x"82007148",x"024002C8",x"CC840000",x"CCA40004",x"CCC40008",x"022002C8",x"C05C0000",x"C0440018",x"8200161C",x"C0620000",x"028002D4",x"C0A20020",x"C82A0000",x"CC280000",x"C0A20020",x"C82A0004",x"CC280004",x"C0A20020",x"C82A0008",x"CC280008",x"02A00001",x"826A7710",x"02A00002",x"826A7648",x"02A00003",x"826A74E8",x"02A00004",x"826A71A8",x"C1FDFFFC",x"C8240000",x"C0620014",x"C8460000",x"44224000",x"C0620010",x"C8460000",x"C49C0000",x"C43C0004",x"C45C0008",x"CC3C0010",x"C17DFFFC",x"40204000",x"03DC0020",x"037E000C",x"C57DFFFC",x"8200083C",x"07DC0020",x"C85C0010",x"48242000",x"C03C0008",x"C8420008",x"C05C0004",x"C0640014",x"C8660008",x"44446000",x"C0640010",x"C8660008",x"CC3C0018",x"CC5C0020",x"C17DFFFC",x"40206000",x"03DC0030",x"037E000C",x"C57DFFFC",x"8200083C",x"07DC0030",x"C85C0020",x"48242000",x"C85C0018",x"48644000",x"48822000",x"40668000",x"8E40725C",x"40804000",x"82007260",x"44804000",x"C8A0006C",x"CCBC0028",x"CC7C0030",x"8E8A7310",x"CC3C0038",x"C17DFFFC",x"40204000",x"03DC0048",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0048",x"C85C0038",x"48242000",x"8E2072A0",x"820072A4",x"44202000",x"C8400068",x"48442000",x"C8600064",x"44446000",x"48442000",x"C8600060",x"44446000",x"48442000",x"C860005C",x"40446000",x"48242000",x"C8400058",x"44224000",x"C8400054",x"48224000",x"C8400050",x"CC3C0040",x"C17DFFFC",x"40204000",x"03DC0050",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0050",x"C85C0040",x"48242000",x"82007314",x"C820004C",x"54220000",x"8E027338",x"58420000",x"8A427330",x"06220001",x"58420000",x"82007334",x"40402000",x"8200733C",x"58420000",x"44224000",x"C03C0008",x"C8420004",x"C03C0004",x"C0420014",x"C8640004",x"44446000",x"C0220010",x"C8620004",x"CC3C0048",x"CC5C0050",x"C17DFFFC",x"40206000",x"03DC0060",x"037E000C",x"C57DFFFC",x"8200083C",x"07DC0060",x"C85C0050",x"48242000",x"C85C0030",x"8E40739C",x"40604000",x"820073A0",x"44604000",x"C89C0028",x"8E687448",x"CC3C0058",x"C17DFFFC",x"40204000",x"03DC0068",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0068",x"C85C0058",x"48242000",x"8E2073D8",x"820073DC",x"44202000",x"C8400068",x"48442000",x"C8600064",x"44446000",x"48442000",x"C8600060",x"44446000",x"48442000",x"C860005C",x"40446000",x"48242000",x"C8400058",x"44224000",x"C8400054",x"48224000",x"C8400050",x"CC3C0060",x"C17DFFFC",x"40204000",x"03DC0070",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0070",x"C85C0060",x"48242000",x"8200744C",x"C820004C",x"54220000",x"8E027470",x"58420000",x"8A427468",x"06220001",x"58420000",x"8200746C",x"40402000",x"82007474",x"58420000",x"44224000",x"C8400048",x"C86000A4",x"C89C0048",x"44868000",x"48888000",x"44448000",x"44262000",x"48222000",x"44242000",x"8E2074A4",x"820074A8",x"40200000",x"C8400044",x"48242000",x"C8400040",x"CC3C0068",x"C17DFFFC",x"40204000",x"03DC0078",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0078",x"C85C0068",x"48242000",x"C03C0000",x"CC220008",x"C1FDFFFC",x"C8240000",x"C0620014",x"C8460000",x"44224000",x"C8440008",x"C0220014",x"C8620008",x"44446000",x"48222000",x"48444000",x"40224000",x"C49C0000",x"C17DFFFC",x"03DC0078",x"037E000C",x"C57DFFFC",x"8200083C",x"07DC0078",x"C840003C",x"CC3C0070",x"C17DFFFC",x"40204000",x"03DC0080",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0080",x"C85C0070",x"48242000",x"54220000",x"8E027580",x"58420000",x"8A427578",x"06220001",x"58420000",x"8200757C",x"40402000",x"82007584",x"58420000",x"44224000",x"C8400050",x"48224000",x"C8400098",x"8E2475B8",x"44224000",x"C17DFFFC",x"03DC0080",x"037E000C",x"C57DFFFC",x"82001270",x"07DC0080",x"82007620",x"8E027604",x"C8600090",x"8E6275E4",x"40224000",x"C17DFFFC",x"03DC0080",x"037E000C",x"C57DFFFC",x"82001270",x"07DC0080",x"82007600",x"02200001",x"C17DFFFC",x"03DC0080",x"037E000C",x"C57DFFFC",x"82000B88",x"07DC0080",x"82007620",x"0220FFFF",x"C17DFFFC",x"03DC0080",x"037E000C",x"C57DFFFC",x"82000B88",x"07DC0080",x"48222000",x"C8400044",x"48624000",x"C03C0000",x"CC620004",x"C86000A8",x"44262000",x"48224000",x"CC220008",x"C1FDFFFC",x"C8240004",x"C8400038",x"48224000",x"C8400098",x"C49C0000",x"8E247680",x"44224000",x"C17DFFFC",x"03DC0080",x"037E000C",x"C57DFFFC",x"82000EC4",x"07DC0080",x"820076E8",x"8E0276CC",x"C8600090",x"8E6276AC",x"40224000",x"C17DFFFC",x"03DC0080",x"037E000C",x"C57DFFFC",x"82000EC4",x"07DC0080",x"820076C8",x"02200001",x"C17DFFFC",x"03DC0080",x"037E000C",x"C57DFFFC",x"8200084C",x"07DC0080",x"820076E8",x"0220FFFF",x"C17DFFFC",x"03DC0080",x"037E000C",x"C57DFFFC",x"8200084C",x"07DC0080",x"48222000",x"C8400044",x"48642000",x"C03C0000",x"CC620000",x"C86000A8",x"44262000",x"48242000",x"CC220004",x"C1FDFFFC",x"C8240000",x"C0620014",x"C8460000",x"44224000",x"C8400034",x"48624000",x"54660000",x"8E067748",x"58860000",x"8A867744",x"06660001",x"58660000",x"82007744",x"8200774C",x"58660000",x"C8800030",x"48668000",x"44226000",x"C860003C",x"C8A40008",x"C0220014",x"C8C20008",x"44AAC000",x"484A4000",x"54240000",x"8E047790",x"58C20000",x"8AC4778C",x"06220001",x"58420000",x"8200778C",x"82007794",x"58420000",x"48448000",x"444A4000",x"8E2677B4",x"8E4677AC",x"C8200044",x"820077B0",x"40200000",x"820077C4",x"8E4677C0",x"40200000",x"820077C4",x"C8200044",x"CC280004",x"C1FDFFFC",x"8E0277D4",x"82007818",x"022002EC",x"024002D4",x"C8820000",x"C8A40000",x"48A2A000",x"4088A000",x"CC820000",x"C8820004",x"C8A40004",x"48A2A000",x"4088A000",x"CC820004",x"C8820008",x"C8A40008",x"4822A000",x"40282000",x"CC220008",x"8E047820",x"C1FDFFFC",x"48244000",x"48222000",x"48226000",x"022002EC",x"C8420000",x"40442000",x"CC420000",x"C8420004",x"40442000",x"CC420004",x"C8420008",x"40242000",x"CC220008",x"C1FDFFFC",x"86207A10",x"02600370",x"22820220",x"D0668000",x"C0860004",x"02A002B4",x"C860002C",x"CC6A0000",x"02C00000",x"02E002A8",x"C10E0000",x"C43C0000",x"CC5C0008",x"C45C0010",x"CC3C0018",x"C49C0020",x"C4FC0024",x"C47C0028",x"C4BC002C",x"C17DFFFC",x"00680000",x"00500000",x"002C0000",x"03DC0038",x"037E000C",x"C57DFFFC",x"820069E8",x"07DC0038",x"C03C002C",x"C8220000",x"C8400070",x"8E4278E0",x"02200000",x"820078F4",x"C8400028",x"8E2478F0",x"02200000",x"820078F4",x"02200001",x"822079F8",x"022002C4",x"C0220000",x"22220220",x"024002B0",x"C0440000",x"00224000",x"C05C0028",x"C0640000",x"82267920",x"820079F4",x"02200000",x"C07C0024",x"C0660000",x"C17DFFFC",x"00460000",x"03DC0038",x"037E000C",x"C57DFFFC",x"82005414",x"07DC0038",x"82207950",x"820079F4",x"022002C8",x"C05C0020",x"C0640000",x"C8220000",x"C8460000",x"48224000",x"C8420004",x"C8660004",x"48446000",x"40224000",x"C8420008",x"C8660008",x"48446000",x"40224000",x"C03C0028",x"C8420008",x"C87C0018",x"48846000",x"48282000",x"C0240000",x"C05C0010",x"C8840000",x"C8A20000",x"4888A000",x"C8A40004",x"C8C20004",x"48AAC000",x"4088A000",x"C8A40008",x"C8C20008",x"48AAC000",x"4088A000",x"48448000",x"C89C0008",x"C17DFFFC",x"40608000",x"03DC0038",x"037E000C",x"C57DFFFC",x"820077CC",x"07DC0038",x"820079F8",x"C03C0000",x"06220001",x"C83C0018",x"C85C0008",x"C05C0010",x"82007858",x"C1FDFFFC",x"02800004",x"86828030",x"C0860008",x"02A002B4",x"C860002C",x"CC6A0000",x"02C00000",x"02E002A8",x"C10E0000",x"CC5C0000",x"C4FC0008",x"C47C000C",x"CC3C0010",x"C45C0018",x"C49C001C",x"C43C0020",x"C4BC0024",x"C17DFFFC",x"00640000",x"002C0000",x"00500000",x"03DC0030",x"037E000C",x"C57DFFFC",x"82005E4C",x"07DC0030",x"C03C0024",x"C8220000",x"C8400070",x"8E427A94",x"02400000",x"82007AA8",x"C8400028",x"8E247AA4",x"02400000",x"82007AA8",x"02400001",x"82407F8C",x"024002C4",x"C0440000",x"026000C8",x"22840220",x"D0668000",x"C0860008",x"C0A6001C",x"C82A0000",x"C85C0010",x"48224000",x"C0A60004",x"02C00001",x"C49C0028",x"CC3C0030",x"C45C0038",x"C47C003C",x"82AC7B50",x"02C00002",x"82AC7B18",x"C17DFFFC",x"00260000",x"03DC0048",x"037E000C",x"C57DFFFC",x"82006F8C",x"07DC0048",x"82007B4C",x"02A002C8",x"C0C60010",x"C86C0000",x"44606000",x"CC6A0000",x"C0C60010",x"C86C0004",x"44606000",x"CC6A0004",x"C0C60010",x"C86C0008",x"44606000",x"CC6A0008",x"82007BA4",x"02A002B0",x"C0AA0000",x"02C002C8",x"CC0C0000",x"CC0C0004",x"CC0C0008",x"06EA0001",x"06AA0001",x"22AA0220",x"C11C0018",x"D870A000",x"8A607B94",x"8E067B8C",x"C860007C",x"82007B90",x"C86000A8",x"82007B98",x"40600000",x"44606000",x"22AE0220",x"DC6CA000",x"0220030C",x"024002B8",x"C8240000",x"CC220000",x"C8240004",x"CC220004",x"C8240008",x"CC220008",x"C03C003C",x"C45C0040",x"C17DFFFC",x"03DC004C",x"037E000C",x"C57DFFFC",x"82007158",x"07DC004C",x"C03C0038",x"22220220",x"024002B0",x"C0440000",x"00224000",x"C05C0020",x"22640220",x"C09C001C",x"D4286000",x"C03C000C",x"C0620004",x"22A40220",x"D066A000",x"C0BC0040",x"C82A0000",x"CC260000",x"C82A0004",x"CC260004",x"C82A0008",x"CC260008",x"C062000C",x"C0DC003C",x"C0EC001C",x"C82E0000",x"C84000A4",x"8E247D0C",x"02E00001",x"23040220",x"D4E70000",x"C0620010",x"22E40220",x"D0E6E000",x"030002D4",x"C8300000",x"CC2E0000",x"C8300004",x"CC2E0004",x"C8300008",x"CC2E0008",x"22E40220",x"D066E000",x"C8200024",x"C47C0044",x"C17DFFFC",x"03DC0050",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0050",x"C85C0030",x"48224000",x"C03C0044",x"C8620000",x"48662000",x"CC620000",x"C8620004",x"48662000",x"CC620004",x"C8620008",x"48262000",x"CC220008",x"C03C000C",x"C042001C",x"C07C0020",x"22860220",x"D0448000",x"028002C8",x"C8280000",x"CC240000",x"C8280004",x"CC240004",x"C8280008",x"CC240008",x"82007D18",x"02E00000",x"23040220",x"D4E70000",x"C8200020",x"024002C8",x"C07C0018",x"C8460000",x"C8640000",x"48446000",x"C8660004",x"C8840004",x"48668000",x"40446000",x"C8660008",x"C8840008",x"48668000",x"40446000",x"48224000",x"C8460000",x"C8640000",x"48626000",x"40446000",x"CC460000",x"C8460004",x"C8640004",x"48626000",x"40446000",x"CC460004",x"C8460008",x"C8640008",x"48226000",x"40242000",x"CC260008",x"C09C003C",x"C0A8001C",x"C82A0004",x"C85C0010",x"48242000",x"02A00000",x"C0DC0008",x"C0CC0000",x"CC3C0048",x"C45C0050",x"C17DFFFC",x"004C0000",x"002A0000",x"03DC005C",x"037E000C",x"C57DFFFC",x"82005414",x"07DC005C",x"82207DE0",x"82007E78",x"022001D0",x"C05C0050",x"C8240000",x"C8420000",x"48224000",x"C8440004",x"C8620004",x"48446000",x"40224000",x"C8440008",x"C8620008",x"48446000",x"40224000",x"44202000",x"C85C0030",x"48224000",x"C05C0018",x"C8640000",x"C8820000",x"48668000",x"C8840004",x"C8A20004",x"4888A000",x"40668000",x"C8840008",x"C8A20008",x"4888A000",x"40668000",x"44606000",x"C89C0048",x"C17DFFFC",x"40406000",x"40608000",x"03DC005C",x"037E000C",x"C57DFFFC",x"820077CC",x"07DC005C",x"02200318",x"C05C0040",x"C8240000",x"CC220000",x"C8240004",x"CC220004",x"C8240008",x"CC220008",x"022000C4",x"C0220000",x"06220001",x"C17DFFFC",x"01240000",x"00420000",x"00320000",x"03DC005C",x"037E000C",x"C57DFFFC",x"8200462C",x"07DC005C",x"02200640",x"C0220000",x"06220001",x"C83C0030",x"C85C0048",x"C05C0018",x"C17DFFFC",x"03DC005C",x"037E000C",x"C57DFFFC",x"82007858",x"07DC005C",x"C820001C",x"C85C0010",x"8E247F08",x"C1FDFFFC",x"02200004",x"C05C0020",x"86427F18",x"82007F2C",x"02240001",x"0260FFFF",x"22220220",x"C09C001C",x"D4682000",x"02200002",x"C07C0028",x"82627F3C",x"82007F88",x"C82000A8",x"C03C003C",x"C022001C",x"C8620000",x"44226000",x"48242000",x"02240001",x"C05C0024",x"C8440000",x"C87C0000",x"40464000",x"C05C0018",x"C07C000C",x"C17DFFFC",x"03DC005C",x"037E000C",x"C57DFFFC",x"82007A14",x"07DC005C",x"C1FDFFFC",x"0220FFFF",x"C05C0020",x"22640220",x"C09C001C",x"D4286000",x"8240802C",x"022001D0",x"C05C0018",x"C8240000",x"C8420000",x"48224000",x"C8440004",x"C8620004",x"48446000",x"40224000",x"C8440008",x"C8620008",x"48446000",x"40224000",x"44202000",x"8E027FE4",x"C1FDFFFC",x"48422000",x"48242000",x"C85C0010",x"48224000",x"022001DC",x"C8420000",x"48224000",x"022002EC",x"C8420000",x"40442000",x"CC420000",x"C8420004",x"40442000",x"CC420004",x"C8420008",x"40242000",x"CC220008",x"C1FDFFFC",x"C1FDFFFC",x"C1FDFFFC",x"024002B4",x"C840002C",x"CC440000",x"02600000",x"028002A8",x"C0A80000",x"CC3C0000",x"C49C0008",x"C43C000C",x"C45C0010",x"C17DFFFC",x"004A0000",x"01260000",x"00620000",x"00320000",x"03DC001C",x"037E000C",x"C57DFFFC",x"820069E8",x"07DC001C",x"C03C0010",x"C8220000",x"C8400070",x"8E42809C",x"02200000",x"820080B0",x"C8400028",x"8E2480AC",x"02200000",x"820080B0",x"02200001",x"8220827C",x"022000C8",x"024002C4",x"C0440000",x"22440220",x"D0224000",x"C05C000C",x"C0440000",x"C0620004",x"02800001",x"C43C0014",x"8268813C",x"02400002",x"82648104",x"C17DFFFC",x"03DC0020",x"037E000C",x"C57DFFFC",x"82006F8C",x"07DC0020",x"82008138",x"024002C8",x"C0620010",x"C8260000",x"44202000",x"CC240000",x"C0620010",x"C8260004",x"44202000",x"CC240004",x"C0620010",x"C8260008",x"44202000",x"CC240008",x"8200818C",x"026002B0",x"C0660000",x"028002C8",x"CC080000",x"CC080004",x"CC080008",x"06A60001",x"06660001",x"22660220",x"D8246000",x"8A20817C",x"8E028174",x"C820007C",x"82008178",x"C82000A8",x"82008180",x"40200000",x"44202000",x"224A0220",x"DC284000",x"024002B8",x"C03C0014",x"C17DFFFC",x"03DC0020",x"037E000C",x"C57DFFFC",x"82007158",x"07DC0020",x"02200000",x"C05C0008",x"C0440000",x"C17DFFFC",x"03DC0020",x"037E000C",x"C57DFFFC",x"82005414",x"07DC0020",x"822081D8",x"C1FDFFFC",x"022002C8",x"024001D0",x"C8220000",x"C8440000",x"48224000",x"C8420004",x"C8640004",x"48446000",x"40224000",x"C8420008",x"C8640008",x"48446000",x"40224000",x"44202000",x"8E02821C",x"40200000",x"8200821C",x"022002E0",x"C85C0000",x"48242000",x"C05C0014",x"C044001C",x"C8440000",x"48224000",x"024002D4",x"C8420000",x"C8640000",x"48626000",x"40446000",x"CC420000",x"C8420004",x"C8640004",x"48626000",x"40446000",x"CC420004",x"C8420008",x"C8640008",x"48226000",x"40242000",x"CC220008",x"C1FDFFFC",x"C1FDFFFC",x"86808490",x"22A80220",x"D0A2A000",x"C0CA0000",x"C82C0000",x"C8440000",x"48224000",x"C84C0004",x"C8640004",x"48446000",x"40224000",x"C84C0008",x"C8640008",x"48446000",x"40224000",x"C47C0000",x"C45C0004",x"C43C0008",x"C49C000C",x"8E208320",x"C8400018",x"C4BC0010",x"CC3C0018",x"C17DFFFC",x"40204000",x"03DC0028",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0028",x"C85C0018",x"48242000",x"C03C0010",x"C17DFFFC",x"03DC0028",x"037E000C",x"C57DFFFC",x"82008034",x"07DC0028",x"82008378",x"02A80001",x"22AA0220",x"D0A2A000",x"C8400014",x"C4BC0020",x"CC3C0018",x"C17DFFFC",x"40204000",x"03DC002C",x"037E000C",x"C57DFFFC",x"82000844",x"07DC002C",x"C85C0018",x"48242000",x"C03C0020",x"C17DFFFC",x"03DC002C",x"037E000C",x"C57DFFFC",x"82008034",x"07DC002C",x"C03C000C",x"06220002",x"8620848C",x"22420220",x"C07C0008",x"D0464000",x"C0840000",x"C8280000",x"C0BC0004",x"C84A0000",x"48224000",x"C8480004",x"C86A0004",x"48446000",x"40224000",x"C8480008",x"C86A0008",x"48446000",x"40224000",x"C43C0024",x"8E20841C",x"C8400018",x"C45C0028",x"CC3C0030",x"C17DFFFC",x"40204000",x"03DC0040",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0040",x"C85C0030",x"48242000",x"C03C0028",x"C17DFFFC",x"03DC0040",x"037E000C",x"C57DFFFC",x"82008034",x"07DC0040",x"82008474",x"02420001",x"22440220",x"D0464000",x"C8400014",x"C45C0038",x"CC3C0030",x"C17DFFFC",x"40204000",x"03DC0044",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0044",x"C85C0030",x"48242000",x"C03C0038",x"C17DFFFC",x"03DC0044",x"037E000C",x"C57DFFFC",x"82008034",x"07DC0044",x"C03C0024",x"06820002",x"C03C0008",x"C05C0004",x"C07C0000",x"82008280",x"C1FDFFFC",x"C1FDFFFC",x"C45C0000",x"C47C0004",x"C43C0008",x"82208524",x"02800354",x"C0880000",x"02A00318",x"C8260000",x"CC2A0000",x"C8260004",x"CC2A0004",x"C8260008",x"CC2A0008",x"02A000C4",x"C0AA0000",x"06AA0001",x"C49C000C",x"C17DFFFC",x"004A0000",x"00260000",x"03DC0018",x"037E000C",x"C57DFFFC",x"8200462C",x"07DC0018",x"02800076",x"C03C000C",x"C05C0000",x"C07C0004",x"C17DFFFC",x"03DC0018",x"037E000C",x"C57DFFFC",x"82008280",x"07DC0018",x"82008524",x"02200001",x"C05C0008",x"824285B4",x"02200354",x"C0220004",x"02600318",x"C09C0004",x"C8280000",x"CC260000",x"C8280004",x"CC260004",x"C8280008",x"CC260008",x"026000C4",x"C0660000",x"06660001",x"C43C0010",x"C17DFFFC",x"00460000",x"00280000",x"03DC001C",x"037E000C",x"C57DFFFC",x"8200462C",x"07DC001C",x"02800076",x"C03C0010",x"C05C0000",x"C07C0004",x"C17DFFFC",x"03DC001C",x"037E000C",x"C57DFFFC",x"82008280",x"07DC001C",x"820085B4",x"02200002",x"C05C0008",x"82428644",x"02200354",x"C0220008",x"02600318",x"C09C0004",x"C8280000",x"CC260000",x"C8280004",x"CC260004",x"C8280008",x"CC260008",x"026000C4",x"C0660000",x"06660001",x"C43C0014",x"C17DFFFC",x"00460000",x"00280000",x"03DC0020",x"037E000C",x"C57DFFFC",x"8200462C",x"07DC0020",x"02800076",x"C03C0014",x"C05C0000",x"C07C0004",x"C17DFFFC",x"03DC0020",x"037E000C",x"C57DFFFC",x"82008280",x"07DC0020",x"82008644",x"02200003",x"C05C0008",x"824286D4",x"02200354",x"C022000C",x"02600318",x"C09C0004",x"C8280000",x"CC260000",x"C8280004",x"CC260004",x"C8280008",x"CC260008",x"026000C4",x"C0660000",x"06660001",x"C43C0018",x"C17DFFFC",x"00460000",x"00280000",x"03DC0024",x"037E000C",x"C57DFFFC",x"8200462C",x"07DC0024",x"02800076",x"C03C0018",x"C05C0000",x"C07C0004",x"C17DFFFC",x"03DC0024",x"037E000C",x"C57DFFFC",x"82008280",x"07DC0024",x"820086D4",x"02200004",x"C05C0008",x"82428748",x"02200354",x"C0220010",x"02400318",x"C07C0004",x"C8260000",x"CC240000",x"C8260004",x"CC240004",x"C8260008",x"CC240008",x"024000C4",x"C0440000",x"06440001",x"C43C001C",x"C17DFFFC",x"00260000",x"03DC0028",x"037E000C",x"C57DFFFC",x"8200462C",x"07DC0028",x"02800076",x"C03C001C",x"C05C0000",x"C07C0004",x"82008280",x"C1FDFFFC",x"C0620014",x"C082001C",x"C0A20004",x"C0C20010",x"02E002E0",x"23040220",x"D0670000",x"C8260000",x"CC2E0000",x"C8260004",x"CC2E0004",x"C8260008",x"CC2E0008",x"C0220018",x"C0220000",x"22640220",x"D0686000",x"22840220",x"D08A8000",x"C4FC0000",x"C4DC0004",x"C45C0008",x"C47C000C",x"C49C0010",x"C43C0014",x"82208914",x"02A00354",x"C0AA0000",x"03000318",x"C8280000",x"CC300000",x"C8280004",x"CC300004",x"C8280008",x"CC300008",x"030000C4",x"C1100000",x"07100001",x"C4BC0018",x"C17DFFFC",x"00500000",x"00280000",x"03DC0024",x"037E000C",x"C57DFFFC",x"8200462C",x"07DC0024",x"C03C0018",x"C04201D8",x"C0640000",x"C8260000",x"C09C000C",x"C8480000",x"48224000",x"C8460004",x"C8680004",x"48446000",x"40224000",x"C8460008",x"C8680008",x"48446000",x"40224000",x"8E208898",x"C8400018",x"C45C001C",x"CC3C0020",x"C17DFFFC",x"40204000",x"03DC0030",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0030",x"C85C0020",x"48242000",x"C03C001C",x"C17DFFFC",x"03DC0030",x"037E000C",x"C57DFFFC",x"82008034",x"07DC0030",x"820088E8",x"C04201DC",x"C8400014",x"C45C0028",x"CC3C0020",x"C17DFFFC",x"40204000",x"03DC0034",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0034",x"C85C0020",x"48242000",x"C03C0028",x"C17DFFFC",x"03DC0034",x"037E000C",x"C57DFFFC",x"82008034",x"07DC0034",x"02800074",x"C03C0018",x"C05C000C",x"C07C0010",x"C17DFFFC",x"03DC0034",x"037E000C",x"C57DFFFC",x"82008280",x"07DC0034",x"82008914",x"02200001",x"C05C0014",x"82428A84",x"02200354",x"C0220004",x"02600318",x"C09C0010",x"C8280000",x"CC260000",x"C8280004",x"CC260004",x"C8280008",x"CC260008",x"026000C4",x"C0660000",x"06660001",x"C43C002C",x"C17DFFFC",x"00460000",x"00280000",x"03DC0038",x"037E000C",x"C57DFFFC",x"8200462C",x"07DC0038",x"C03C002C",x"C04201D8",x"C0640000",x"C8260000",x"C09C000C",x"C8480000",x"48224000",x"C8460004",x"C8680004",x"48446000",x"40224000",x"C8460008",x"C8680008",x"48446000",x"40224000",x"8E208A08",x"C8400018",x"C45C0030",x"CC3C0038",x"C17DFFFC",x"40204000",x"03DC0048",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0048",x"C85C0038",x"48242000",x"C03C0030",x"C17DFFFC",x"03DC0048",x"037E000C",x"C57DFFFC",x"82008034",x"07DC0048",x"82008A58",x"C04201DC",x"C8400014",x"C45C0040",x"CC3C0038",x"C17DFFFC",x"40204000",x"03DC004C",x"037E000C",x"C57DFFFC",x"82000844",x"07DC004C",x"C85C0038",x"48242000",x"C03C0040",x"C17DFFFC",x"03DC004C",x"037E000C",x"C57DFFFC",x"82008034",x"07DC004C",x"02800074",x"C03C002C",x"C05C000C",x"C07C0010",x"C17DFFFC",x"03DC004C",x"037E000C",x"C57DFFFC",x"82008280",x"07DC004C",x"82008A84",x"02200002",x"C05C0014",x"82428BF4",x"02200354",x"C0220008",x"02600318",x"C09C0010",x"C8280000",x"CC260000",x"C8280004",x"CC260004",x"C8280008",x"CC260008",x"026000C4",x"C0660000",x"06660001",x"C43C0044",x"C17DFFFC",x"00460000",x"00280000",x"03DC0050",x"037E000C",x"C57DFFFC",x"8200462C",x"07DC0050",x"C03C0044",x"C04201D8",x"C0640000",x"C8260000",x"C09C000C",x"C8480000",x"48224000",x"C8460004",x"C8680004",x"48446000",x"40224000",x"C8460008",x"C8680008",x"48446000",x"40224000",x"8E208B78",x"C8400018",x"C45C0048",x"CC3C0050",x"C17DFFFC",x"40204000",x"03DC0060",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0060",x"C85C0050",x"48242000",x"C03C0048",x"C17DFFFC",x"03DC0060",x"037E000C",x"C57DFFFC",x"82008034",x"07DC0060",x"82008BC8",x"C04201DC",x"C8400014",x"C45C0058",x"CC3C0050",x"C17DFFFC",x"40204000",x"03DC0064",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0064",x"C85C0050",x"48242000",x"C03C0058",x"C17DFFFC",x"03DC0064",x"037E000C",x"C57DFFFC",x"82008034",x"07DC0064",x"02800074",x"C03C0044",x"C05C000C",x"C07C0010",x"C17DFFFC",x"03DC0064",x"037E000C",x"C57DFFFC",x"82008280",x"07DC0064",x"82008BF4",x"02200003",x"C05C0014",x"82428D64",x"02200354",x"C022000C",x"02600318",x"C09C0010",x"C8280000",x"CC260000",x"C8280004",x"CC260004",x"C8280008",x"CC260008",x"026000C4",x"C0660000",x"06660001",x"C43C005C",x"C17DFFFC",x"00460000",x"00280000",x"03DC0068",x"037E000C",x"C57DFFFC",x"8200462C",x"07DC0068",x"C03C005C",x"C04201D8",x"C0640000",x"C8260000",x"C09C000C",x"C8480000",x"48224000",x"C8460004",x"C8680004",x"48446000",x"40224000",x"C8460008",x"C8680008",x"48446000",x"40224000",x"8E208CE8",x"C8400018",x"C45C0060",x"CC3C0068",x"C17DFFFC",x"40204000",x"03DC0078",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0078",x"C85C0068",x"48242000",x"C03C0060",x"C17DFFFC",x"03DC0078",x"037E000C",x"C57DFFFC",x"82008034",x"07DC0078",x"82008D38",x"C04201DC",x"C8400014",x"C45C0070",x"CC3C0068",x"C17DFFFC",x"40204000",x"03DC007C",x"037E000C",x"C57DFFFC",x"82000844",x"07DC007C",x"C85C0068",x"48242000",x"C03C0070",x"C17DFFFC",x"03DC007C",x"037E000C",x"C57DFFFC",x"82008034",x"07DC007C",x"02800074",x"C03C005C",x"C05C000C",x"C07C0010",x"C17DFFFC",x"03DC007C",x"037E000C",x"C57DFFFC",x"82008280",x"07DC007C",x"82008D64",x"02200004",x"C05C0014",x"82428ED0",x"02200354",x"C0220010",x"02400318",x"C07C0010",x"C8260000",x"CC240000",x"C8260004",x"CC240004",x"C8260008",x"CC240008",x"024000C4",x"C0440000",x"06440001",x"C43C0074",x"C17DFFFC",x"00260000",x"03DC0080",x"037E000C",x"C57DFFFC",x"8200462C",x"07DC0080",x"C03C0074",x"C04201D8",x"C0640000",x"C8260000",x"C09C000C",x"C8480000",x"48224000",x"C8460004",x"C8680004",x"48446000",x"40224000",x"C8460008",x"C8680008",x"48446000",x"40224000",x"8E208E54",x"C8400018",x"C45C0078",x"CC3C0080",x"C17DFFFC",x"40204000",x"03DC0090",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0090",x"C85C0080",x"48242000",x"C03C0078",x"C17DFFFC",x"03DC0090",x"037E000C",x"C57DFFFC",x"82008034",x"07DC0090",x"82008EA4",x"C04201DC",x"C8400014",x"C45C0088",x"CC3C0080",x"C17DFFFC",x"40204000",x"03DC0094",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0094",x"C85C0080",x"48242000",x"C03C0088",x"C17DFFFC",x"03DC0094",x"037E000C",x"C57DFFFC",x"82008034",x"07DC0094",x"02800074",x"C03C0074",x"C05C000C",x"C07C0010",x"C17DFFFC",x"03DC0094",x"037E000C",x"C57DFFFC",x"82008280",x"07DC0094",x"82008ED0",x"022002EC",x"C05C0008",x"22440220",x"C07C0004",x"D0464000",x"C8220000",x"C8440000",x"C07C0000",x"C8660000",x"48446000",x"40224000",x"CC220000",x"C8220004",x"C8440004",x"C8660004",x"48446000",x"40224000",x"CC220004",x"C8220008",x"C8440008",x"C8660008",x"48446000",x"40224000",x"CC220008",x"C1FDFFFC",x"22C20220",x"D044C000",x"C0440014",x"06C20001",x"22CC0220",x"D0C6C000",x"C0CC0014",x"22E20220",x"D0E6E000",x"C0EE0014",x"03020001",x"23100220",x"D1070000",x"C1100014",x"23220220",x"D0892000",x"C0880014",x"032002E0",x"234A0220",x"D0454000",x"C8240000",x"CC320000",x"C8240004",x"CC320004",x"C8240008",x"CC320008",x"224A0220",x"D04C4000",x"C8320000",x"C8440000",x"40224000",x"CC320000",x"C8320004",x"C8440004",x"40224000",x"CC320004",x"C8320008",x"C8440008",x"40224000",x"CC320008",x"224A0220",x"D04E4000",x"C8320000",x"C8440000",x"40224000",x"CC320000",x"C8320004",x"C8440004",x"40224000",x"CC320004",x"C8320008",x"C8440008",x"40224000",x"CC320008",x"224A0220",x"D0504000",x"C8320000",x"C8440000",x"40224000",x"CC320000",x"C8320004",x"C8440004",x"40224000",x"CC320004",x"C8320008",x"C8440008",x"40224000",x"CC320008",x"224A0220",x"D0484000",x"C8320000",x"C8440000",x"40224000",x"CC320000",x"C8320004",x"C8440004",x"40224000",x"CC320004",x"C8320008",x"C8440008",x"40224000",x"CC320008",x"22220220",x"D0262000",x"C0220010",x"024002EC",x"226A0220",x"D0226000",x"C8240000",x"C8420000",x"C8720000",x"48446000",x"40224000",x"CC240000",x"C8240004",x"C8420004",x"C8720004",x"48446000",x"40224000",x"CC240004",x"C8240008",x"C8420008",x"C8720008",x"48446000",x"40224000",x"CC240008",x"C1FDFFFC",x"02600004",x"86649258",x"C0620008",x"22840220",x"D0668000",x"86609254",x"C062000C",x"22840220",x"D0668000",x"C43C0000",x"826091EC",x"C0620014",x"C082001C",x"C0A20004",x"C0C20010",x"02E002E0",x"23040220",x"D0670000",x"C8260000",x"CC2E0000",x"C8260004",x"CC2E0004",x"C8260008",x"CC2E0008",x"C0620018",x"C0660000",x"23040220",x"D0890000",x"23040220",x"D0AB0000",x"C4FC0004",x"C4DC0008",x"C45C000C",x"C17DFFFC",x"00480000",x"00260000",x"006A0000",x"03DC0018",x"037E000C",x"C57DFFFC",x"82008494",x"07DC0018",x"022002EC",x"C05C000C",x"22640220",x"C09C0008",x"D0686000",x"C8220000",x"C8460000",x"C09C0004",x"C8680000",x"48446000",x"40224000",x"CC220000",x"C8220004",x"C8460004",x"C8680004",x"48446000",x"40224000",x"CC220004",x"C8220008",x"C8460008",x"C8680008",x"48446000",x"40224000",x"CC220008",x"820091EC",x"02440001",x"02200004",x"86249250",x"C03C0000",x"C0620008",x"22840220",x"D0668000",x"8660924C",x"C062000C",x"22840220",x"D0668000",x"C45C0010",x"8260923C",x"C17DFFFC",x"03DC001C",x"037E000C",x"C57DFFFC",x"8200874C",x"07DC001C",x"8200923C",x"C03C0010",x"02420001",x"C03C0000",x"820090E0",x"C1FDFFFC",x"C1FDFFFC",x"C1FDFFFC",x"C1FDFFFC",x"22E20220",x"D0E8E000",x"03000004",x"870C9528",x"C10E0008",x"232C0220",x"D1112000",x"87009524",x"C10E0008",x"232C0220",x"D1112000",x"23220220",x"D1272000",x"C1320008",x"234C0220",x"D1334000",x"833092A8",x"03000000",x"82009314",x"23220220",x"D12B2000",x"C1320008",x"234C0220",x"D1334000",x"833092C8",x"03000000",x"82009314",x"07220001",x"23320220",x"D1292000",x"C1320008",x"234C0220",x"D1334000",x"833092EC",x"03000000",x"82009314",x"03220001",x"23320220",x"D1292000",x"C1320008",x"234C0220",x"D1334000",x"83309310",x"03000000",x"82009314",x"03000001",x"830094B8",x"C0EE000C",x"230C0220",x"D0EF0000",x"C45C0000",x"C4BC0004",x"C47C0008",x"C49C000C",x"C43C0010",x"C4DC0014",x"82E0936C",x"C17DFFFC",x"00460000",x"00680000",x"008A0000",x"00AC0000",x"03DC0020",x"037E000C",x"C57DFFFC",x"82008F34",x"07DC0020",x"8200936C",x"C03C0014",x"02420001",x"C03C0010",x"22620220",x"C09C000C",x"D0686000",x"02A00004",x"86A494B4",x"C0A60008",x"22C40220",x"D0AAC000",x"86A094B0",x"C0A60008",x"22C40220",x"D0AAC000",x"22C20220",x"C0FC0008",x"D0CEC000",x"C0CC0008",x"23040220",x"D0CD0000",x"82CA93CC",x"02A00000",x"8200943C",x"22C20220",x"C11C0004",x"D0D0C000",x"C0CC0008",x"23240220",x"D0CD2000",x"82CA93F0",x"02A00000",x"8200943C",x"06C20001",x"22CC0220",x"D0C8C000",x"C0CC0008",x"23240220",x"D0CD2000",x"82CA9414",x"02A00000",x"8200943C",x"02C20001",x"22CC0220",x"D0C8C000",x"C0CC0008",x"23240220",x"D0CD2000",x"82CA9438",x"02A00000",x"8200943C",x"02A00001",x"82A094A8",x"C066000C",x"22A40220",x"D066A000",x"C45C0018",x"82609488",x"C07C0004",x"C17DFFFC",x"00A40000",x"004E0000",x"01280000",x"00860000",x"00720000",x"03DC0024",x"037E000C",x"C57DFFFC",x"82008F34",x"07DC0024",x"82009488",x"C03C0018",x"02C20001",x"C03C0010",x"C05C0000",x"C07C0008",x"C09C000C",x"C0BC0004",x"8200925C",x"00260000",x"820090E0",x"C1FDFFFC",x"C1FDFFFC",x"02200004",x"862C9520",x"C02E0008",x"224C0220",x"D0224000",x"8620951C",x"C02E000C",x"224C0220",x"D0224000",x"C4FC001C",x"C4DC0014",x"8220950C",x"C17DFFFC",x"004C0000",x"002E0000",x"03DC0028",x"037E000C",x"C57DFFFC",x"8200874C",x"07DC0028",x"8200950C",x"C03C0014",x"02420001",x"C03C001C",x"820090E0",x"C1FDFFFC",x"C1FDFFFC",x"C1FDFFFC",x"C1FDFFFC",x"02600004",x"8664986C",x"C0620008",x"22840220",x"D0668000",x"86609868",x"C062000C",x"22840220",x"D0668000",x"C45C0000",x"8260964C",x"C0620018",x"C0660000",x"028002E0",x"CC080000",x"CC080004",x"CC080008",x"C0A2001C",x"C0C20004",x"02E00354",x"22660220",x"D06E6000",x"22E40220",x"D0AAE000",x"22E40220",x"D0CCE000",x"02E00318",x"C82C0000",x"CC2E0000",x"C82C0004",x"CC2E0004",x"C82C0008",x"CC2E0008",x"02E000C4",x"C0EE0000",x"06EE0001",x"C49C0004",x"C43C0008",x"C4DC000C",x"C4BC0010",x"C47C0014",x"C17DFFFC",x"004E0000",x"002C0000",x"03DC0020",x"037E000C",x"C57DFFFC",x"8200462C",x"07DC0020",x"02800076",x"C03C0014",x"C05C0010",x"C07C000C",x"C17DFFFC",x"03DC0020",x"037E000C",x"C57DFFFC",x"82008280",x"07DC0020",x"C03C0008",x"C0420014",x"C07C0000",x"22860220",x"D0448000",x"C09C0004",x"C8280000",x"CC240000",x"C8280004",x"CC240004",x"C8280008",x"CC240008",x"8200964C",x"C05C0000",x"02440001",x"02600004",x"86649864",x"C0620008",x"22840220",x"D0668000",x"86609860",x"C062000C",x"22840220",x"D0668000",x"C45C0018",x"82609854",x"C0620018",x"C0660000",x"028002E0",x"CC080000",x"CC080004",x"CC080008",x"C0A2001C",x"C0C20004",x"02E00354",x"22660220",x"D06E6000",x"22E40220",x"D0AAE000",x"22E40220",x"D0CCE000",x"02E00318",x"C82C0000",x"CC2E0000",x"C82C0004",x"CC2E0004",x"C82C0008",x"CC2E0008",x"02E000C4",x"C0EE0000",x"06EE0001",x"C49C001C",x"C43C0008",x"C4DC0020",x"C4BC0024",x"C47C0028",x"C17DFFFC",x"004E0000",x"002C0000",x"03DC0034",x"037E000C",x"C57DFFFC",x"8200462C",x"07DC0034",x"C03C0028",x"C04201D8",x"C0640000",x"C8260000",x"C09C0024",x"C8480000",x"48224000",x"C8460004",x"C8680004",x"48446000",x"40224000",x"C8460008",x"C8680008",x"48446000",x"40224000",x"8E2097A8",x"C8400018",x"C45C002C",x"CC3C0030",x"C17DFFFC",x"40204000",x"03DC0040",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0040",x"C85C0030",x"48242000",x"C03C002C",x"C17DFFFC",x"03DC0040",x"037E000C",x"C57DFFFC",x"82008034",x"07DC0040",x"820097F8",x"C04201DC",x"C8400014",x"C45C0038",x"CC3C0030",x"C17DFFFC",x"40204000",x"03DC0044",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0044",x"C85C0030",x"48242000",x"C03C0038",x"C17DFFFC",x"03DC0044",x"037E000C",x"C57DFFFC",x"82008034",x"07DC0044",x"02800074",x"C03C0028",x"C05C0024",x"C07C0020",x"C17DFFFC",x"03DC0044",x"037E000C",x"C57DFFFC",x"82008280",x"07DC0044",x"C03C0008",x"C0420014",x"C07C0018",x"22860220",x"D0448000",x"C09C001C",x"C8280000",x"CC240000",x"C8280004",x"CC240004",x"C8280008",x"CC240008",x"82009854",x"C05C0018",x"02440001",x"8200952C",x"C1FDFFFC",x"C1FDFFFC",x"C1FDFFFC",x"C1FDFFFC",x"86409C04",x"02800308",x"C8880000",x"02800300",x"C0880000",x"04848000",x"58A80000",x"4888A000",x"02800348",x"02A00324",x"C8AA0000",x"48A8A000",x"40AA2000",x"CCA80000",x"C8AA0004",x"48A8A000",x"40AA4000",x"CCA80004",x"C8AA0008",x"4888A000",x"40886000",x"CC880008",x"02A00000",x"CC7C0000",x"CC5C0008",x"CC3C0010",x"C47C0018",x"C49C001C",x"C43C0020",x"C45C0024",x"C17DFFFC",x"004A0000",x"00280000",x"03DC0030",x"037E000C",x"C57DFFFC",x"8200161C",x"07DC0030",x"022002EC",x"40400000",x"CC020000",x"CC020004",x"CC020008",x"0240030C",x"026001C4",x"C8260000",x"CC240000",x"C8260004",x"CC240004",x"C8260008",x"CC240008",x"02400000",x"C82000A8",x"C07C0024",x"22860220",x"C0BC0020",x"D08A8000",x"C0DC001C",x"C43C0028",x"C17DFFFC",x"00680000",x"00240000",x"004C0000",x"03DC0034",x"037E000C",x"C57DFFFC",x"82007A14",x"07DC0034",x"C03C0024",x"22420220",x"C07C0020",x"D0464000",x"C0440000",x"C09C0028",x"C8280000",x"CC240000",x"C8280004",x"CC240004",x"C8280008",x"CC240008",x"22420220",x"D0464000",x"C0440018",x"C09C0018",x"C4840000",x"22420220",x"D0464000",x"C0A40008",x"C0AA0000",x"86A09BCC",x"C0A4000C",x"C0AA0000",x"C45C002C",x"82A09BA8",x"C0A40018",x"C0AA0000",x"02C002E0",x"CC0C0000",x"CC0C0004",x"CC0C0008",x"C0E4001C",x"C1040004",x"03200354",x"22AA0220",x"D0B2A000",x"C0EE0000",x"C1100000",x"03200318",x"C8300000",x"CC320000",x"C8300004",x"CC320004",x"C8300008",x"CC320008",x"032000C4",x"C1320000",x"07320001",x"C4DC0030",x"C51C0034",x"C4FC0038",x"C4BC003C",x"C17DFFFC",x"00520000",x"00300000",x"03DC0048",x"037E000C",x"C57DFFFC",x"8200462C",x"07DC0048",x"C03C003C",x"C04201D8",x"C0640000",x"C8260000",x"C09C0038",x"C8480000",x"48224000",x"C8460004",x"C8680004",x"48446000",x"40224000",x"C8460008",x"C8680008",x"48446000",x"40224000",x"8E209B04",x"C8400018",x"C45C0040",x"CC3C0048",x"C17DFFFC",x"40204000",x"03DC0058",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0058",x"C85C0048",x"48242000",x"C03C0040",x"C17DFFFC",x"03DC0058",x"037E000C",x"C57DFFFC",x"82008034",x"07DC0058",x"82009B54",x"C04201DC",x"C8400014",x"C45C0050",x"CC3C0048",x"C17DFFFC",x"40204000",x"03DC005C",x"037E000C",x"C57DFFFC",x"82000844",x"07DC005C",x"C85C0048",x"48242000",x"C03C0050",x"C17DFFFC",x"03DC005C",x"037E000C",x"C57DFFFC",x"82008034",x"07DC005C",x"02800074",x"C03C003C",x"C05C0038",x"C07C0034",x"C17DFFFC",x"03DC005C",x"037E000C",x"C57DFFFC",x"82008280",x"07DC005C",x"C03C002C",x"C0420014",x"C0440000",x"C07C0030",x"C8260000",x"CC240000",x"C8260004",x"CC240004",x"C8260008",x"CC240008",x"82009BA8",x"02400001",x"C03C002C",x"C17DFFFC",x"03DC005C",x"037E000C",x"C57DFFFC",x"8200952C",x"07DC005C",x"82009BCC",x"C03C0024",x"06420001",x"C03C0018",x"02220001",x"02600005",x"86269BEC",x"06620005",x"82009BF0",x"00620000",x"C83C0010",x"C85C0008",x"C87C0000",x"C03C0020",x"82009870",x"C1FDFFFC",x"02800308",x"C8280000",x"02800300",x"C0880004",x"04448000",x"58440000",x"48224000",x"02400330",x"C8440000",x"48424000",x"0280033C",x"C8680000",x"40446000",x"C8640004",x"48626000",x"C8880004",x"40668000",x"C8840008",x"48228000",x"C8880008",x"40228000",x"024002F8",x"C0440000",x"06440001",x"41E06000",x"40602000",x"40204000",x"4041E000",x"82009870",x"02C002F8",x"C0EC0000",x"862E9C8C",x"C1FDFFFC",x"02E002EC",x"23020220",x"D1090000",x"C1100000",x"C8300000",x"CC2E0000",x"C8300004",x"CC2E0004",x"C8300008",x"CC2E0008",x"03040001",x"C12C0004",x"87129CC8",x"03000000",x"82009CF8",x"86049CD4",x"03000000",x"82009CF8",x"03020001",x"C12C0000",x"87129CE8",x"03000000",x"82009CF8",x"86029CF4",x"03000000",x"82009CF8",x"03000001",x"C4BC0000",x"C47C0004",x"C45C0008",x"C49C000C",x"C4DC0010",x"C43C0014",x"C4FC0018",x"83009E4C",x"03000000",x"23220220",x"D1292000",x"C1520008",x"C1540000",x"87409E48",x"C1520008",x"C1540000",x"22C20220",x"D0C6C000",x"C0CC0008",x"C0CC0000",x"82D49D54",x"02C00000",x"82009DB4",x"22C20220",x"D0CAC000",x"C0CC0008",x"C0CC0000",x"82D49D70",x"02C00000",x"82009DB4",x"06C20001",x"22CC0220",x"D0C8C000",x"C0CC0008",x"C0CC0000",x"82D49D90",x"02C00000",x"82009DB4",x"02C20001",x"22CC0220",x"D0C8C000",x"C0CC0008",x"C0CC0000",x"82D49DB0",x"02C00000",x"82009DB4",x"02C00001",x"82C09E24",x"C0D2000C",x"C0CC0000",x"82C09DF0",x"C17DFFFC",x"00460000",x"00680000",x"008A0000",x"00B00000",x"03DC0024",x"037E000C",x"C57DFFFC",x"82008F34",x"07DC0024",x"82009DF0",x"02C00001",x"C03C0014",x"C05C0008",x"C07C0004",x"C09C000C",x"C0BC0000",x"C17DFFFC",x"03DC0024",x"037E000C",x"C57DFFFC",x"8200925C",x"07DC0024",x"82009E44",x"C17DFFFC",x"00500000",x"00320000",x"03DC0024",x"037E000C",x"C57DFFFC",x"820090E0",x"07DC0024",x"82009E48",x"82009EBC",x"23020220",x"D1090000",x"03200000",x"C1500008",x"C1540000",x"87409EBC",x"C150000C",x"C1540000",x"C51C001C",x"83409E98",x"C17DFFFC",x"00520000",x"00300000",x"03DC0028",x"037E000C",x"C57DFFFC",x"8200874C",x"07DC0028",x"82009E98",x"02400001",x"C03C001C",x"C17DFFFC",x"03DC0028",x"037E000C",x"C57DFFFC",x"820090E0",x"07DC0028",x"82009EBC",x"C03C0018",x"C8220000",x"54420000",x"026000FF",x"86649EE0",x"86409ED8",x"82009EDC",x"02400000",x"82009EE4",x"024000FF",x"C17DFFFC",x"00240000",x"03DC0028",x"037E000C",x"C57DFFFC",x"8200078C",x"07DC0028",x"C03C0018",x"C8220004",x"54420000",x"026000FF",x"86649F24",x"86409F1C",x"82009F20",x"02400000",x"82009F28",x"024000FF",x"C17DFFFC",x"00240000",x"03DC0028",x"037E000C",x"C57DFFFC",x"8200078C",x"07DC0028",x"C03C0018",x"C8220008",x"54420000",x"026000FF",x"86649F68",x"86409F60",x"82009F64",x"02400000",x"82009F6C",x"024000FF",x"C17DFFFC",x"00240000",x"03DC0028",x"037E000C",x"C57DFFFC",x"8200078C",x"07DC0028",x"C03C0014",x"02220001",x"C05C0010",x"C0640000",x"86269FA0",x"C1FDFFFC",x"22620220",x"C09C000C",x"D0686000",x"C0660000",x"C8260000",x"C0BC0018",x"CC2A0000",x"C8260004",x"CC2A0004",x"C8260008",x"CC2A0008",x"C07C0008",x"02C60001",x"C0E40004",x"86CE9FE4",x"02400000",x"8200A014",x"86069FF0",x"02400000",x"8200A014",x"02C20001",x"C0440000",x"86C4A004",x"02400000",x"8200A014",x"8602A010",x"02400000",x"8200A014",x"02400001",x"C43C0020",x"8240A054",x"02C00000",x"C05C0004",x"C0FC0000",x"C17DFFFC",x"00AE0000",x"01260000",x"00640000",x"00520000",x"03DC002C",x"037E000C",x"C57DFFFC",x"8200925C",x"07DC002C",x"8200A080",x"22420220",x"D0484000",x"02C00000",x"C17DFFFC",x"00240000",x"004C0000",x"03DC002C",x"037E000C",x"C57DFFFC",x"820090E0",x"07DC002C",x"C03C0018",x"C8220000",x"54420000",x"026000FF",x"8664A0A4",x"8640A09C",x"8200A0A0",x"02400000",x"8200A0A8",x"024000FF",x"C17DFFFC",x"00240000",x"03DC002C",x"037E000C",x"C57DFFFC",x"8200078C",x"07DC002C",x"C03C0018",x"C8220004",x"54420000",x"026000FF",x"8664A0E8",x"8640A0E0",x"8200A0E4",x"02400000",x"8200A0EC",x"024000FF",x"C17DFFFC",x"00240000",x"03DC002C",x"037E000C",x"C57DFFFC",x"8200078C",x"07DC002C",x"C03C0018",x"C8220008",x"54220000",x"024000FF",x"8642A12C",x"8620A124",x"8200A128",x"02200000",x"8200A130",x"022000FF",x"C17DFFFC",x"03DC002C",x"037E000C",x"C57DFFFC",x"8200078C",x"07DC002C",x"C03C0020",x"02220001",x"C05C0008",x"C07C0004",x"C09C000C",x"C0BC0000",x"82009C7C",x"02C002F8",x"C0EC0004",x"862EA174",x"C1FDFFFC",x"C0EC0004",x"06EE0001",x"C4BC0000",x"C49C0004",x"C45C0008",x"C43C000C",x"C47C0010",x"C4DC0014",x"862EA19C",x"8200A1C4",x"02E20001",x"C17DFFFC",x"006A0000",x"004E0000",x"00280000",x"03DC0020",x"037E000C",x"C57DFFFC",x"82009C08",x"07DC0020",x"02200000",x"C05C0014",x"C0640000",x"8606A1D8",x"8200A390",x"026002EC",x"C09C0010",x"C0A80000",x"C0AA0000",x"C82A0000",x"CC260000",x"C82A0004",x"CC260004",x"C82A0008",x"CC260008",x"C0BC000C",x"02CA0001",x"C0E40004",x"86CEA218",x"02C00000",x"8200A23C",x"860AA224",x"02C00000",x"8200A23C",x"02C00001",x"C0E40000",x"86CEA238",x"02C00000",x"8200A23C",x"02C00001",x"C47C0018",x"82C0A278",x"02C00000",x"C0FC0008",x"C11C0004",x"C17DFFFC",x"006E0000",x"004A0000",x"00B00000",x"03DC0024",x"037E000C",x"C57DFFFC",x"8200925C",x"07DC0024",x"8200A29C",x"C0280000",x"02C00000",x"C17DFFFC",x"004C0000",x"03DC0024",x"037E000C",x"C57DFFFC",x"820090E0",x"07DC0024",x"C03C0018",x"C8220000",x"54420000",x"026000FF",x"8664A2C0",x"8640A2B8",x"8200A2BC",x"02400000",x"8200A2C4",x"024000FF",x"C17DFFFC",x"00240000",x"03DC0024",x"037E000C",x"C57DFFFC",x"8200078C",x"07DC0024",x"C03C0018",x"C8220004",x"54420000",x"026000FF",x"8664A304",x"8640A2FC",x"8200A300",x"02400000",x"8200A308",x"024000FF",x"C17DFFFC",x"00240000",x"03DC0024",x"037E000C",x"C57DFFFC",x"8200078C",x"07DC0024",x"C03C0018",x"C8220008",x"54220000",x"024000FF",x"8642A348",x"8620A340",x"8200A344",x"02200000",x"8200A34C",x"022000FF",x"C17DFFFC",x"03DC0024",x"037E000C",x"C57DFFFC",x"8200078C",x"07DC0024",x"02200001",x"C05C000C",x"C07C0008",x"C09C0010",x"C0BC0004",x"C17DFFFC",x"03DC0024",x"037E000C",x"C57DFFFC",x"82009C7C",x"07DC0024",x"C03C000C",x"02420001",x"C03C0000",x"02220002",x"02600005",x"8626A3B0",x"06620005",x"8200A3B4",x"00620000",x"C03C0014",x"C0820004",x"8648A3C4",x"8200A478",x"C0220004",x"06220001",x"C47C001C",x"C45C0020",x"8642A3DC",x"8200A404",x"02240001",x"C09C0008",x"C17DFFFC",x"00420000",x"00280000",x"03DC002C",x"037E000C",x"C57DFFFC",x"82009C08",x"07DC002C",x"02200000",x"C05C0020",x"C07C0010",x"C09C0004",x"C0BC0008",x"C17DFFFC",x"03DC002C",x"037E000C",x"C57DFFFC",x"82009C7C",x"07DC002C",x"C03C0020",x"02220001",x"C05C001C",x"02440002",x"02600005",x"8646A450",x"06A40005",x"8200A454",x"00A40000",x"C05C0004",x"C07C0008",x"C09C0010",x"C17DFFFC",x"03DC002C",x"037E000C",x"C57DFFFC",x"8200A164",x"07DC002C",x"C1FDFFFC",x"02200003",x"40200000",x"CC3C0000",x"C17DFFFC",x"03DC0010",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0010",x"02400003",x"C83C0000",x"C43C0008",x"C17DFFFC",x"00240000",x"03DC0014",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0014",x"00420000",x"02200005",x"C17DFFFC",x"03DC0014",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0014",x"02400003",x"C83C0000",x"C43C000C",x"C17DFFFC",x"00240000",x"03DC0018",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0018",x"C05C000C",x"C4240004",x"02200003",x"C83C0000",x"C17DFFFC",x"03DC0018",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0018",x"C05C000C",x"C4240008",x"02200003",x"C83C0000",x"C17DFFFC",x"03DC0018",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0018",x"C05C000C",x"C424000C",x"02200003",x"C83C0000",x"C17DFFFC",x"03DC0018",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0018",x"C05C000C",x"C4240010",x"02200005",x"02600000",x"C17DFFFC",x"00460000",x"03DC0018",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0018",x"02400005",x"02600000",x"C43C0010",x"C17DFFFC",x"00240000",x"00460000",x"03DC001C",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC001C",x"02400003",x"C83C0000",x"C43C0014",x"C17DFFFC",x"00240000",x"03DC0020",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0020",x"00420000",x"02200005",x"C17DFFFC",x"03DC0020",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0020",x"02400003",x"C83C0000",x"C43C0018",x"C17DFFFC",x"00240000",x"03DC0024",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0024",x"C05C0018",x"C4240004",x"02200003",x"C83C0000",x"C17DFFFC",x"03DC0024",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0024",x"C05C0018",x"C4240008",x"02200003",x"C83C0000",x"C17DFFFC",x"03DC0024",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0024",x"C05C0018",x"C424000C",x"02200003",x"C83C0000",x"C17DFFFC",x"03DC0024",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0024",x"C05C0018",x"C4240010",x"02200003",x"C83C0000",x"C17DFFFC",x"03DC0024",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0024",x"00420000",x"02200005",x"C17DFFFC",x"03DC0024",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0024",x"02400003",x"C83C0000",x"C43C001C",x"C17DFFFC",x"00240000",x"03DC0028",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0028",x"C05C001C",x"C4240004",x"02200003",x"C83C0000",x"C17DFFFC",x"03DC0028",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0028",x"C05C001C",x"C4240008",x"02200003",x"C83C0000",x"C17DFFFC",x"03DC0028",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0028",x"C05C001C",x"C424000C",x"02200003",x"C83C0000",x"C17DFFFC",x"03DC0028",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0028",x"C05C001C",x"C4240010",x"02200001",x"02600000",x"C17DFFFC",x"00460000",x"03DC0028",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0028",x"02400003",x"C83C0000",x"C43C0020",x"C17DFFFC",x"00240000",x"03DC002C",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC002C",x"00420000",x"02200005",x"C17DFFFC",x"03DC002C",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC002C",x"02400003",x"C83C0000",x"C43C0024",x"C17DFFFC",x"00240000",x"03DC0030",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0030",x"C05C0024",x"C4240004",x"02200003",x"C83C0000",x"C17DFFFC",x"03DC0030",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0030",x"C05C0024",x"C4240008",x"02200003",x"C83C0000",x"C17DFFFC",x"03DC0030",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0030",x"C05C0024",x"C424000C",x"02200003",x"C83C0000",x"C17DFFFC",x"03DC0030",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0030",x"C05C0024",x"C4240010",x"003A0000",x"03BA0020",x"C442001C",x"C05C0020",x"C4420018",x"C05C001C",x"C4420014",x"C05C0018",x"C4420010",x"C05C0014",x"C442000C",x"C05C0010",x"C4420008",x"C05C000C",x"C4420004",x"C05C0008",x"C4420000",x"C1FDFFFC",x"8640AE10",x"02600003",x"40200000",x"C43C0000",x"C45C0004",x"CC3C0008",x"C17DFFFC",x"00260000",x"03DC0018",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0018",x"02400003",x"C83C0008",x"C43C0010",x"C17DFFFC",x"00240000",x"03DC001C",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC001C",x"00420000",x"02200005",x"C17DFFFC",x"03DC001C",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC001C",x"02400003",x"C83C0008",x"C43C0014",x"C17DFFFC",x"00240000",x"03DC0020",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0020",x"C05C0014",x"C4240004",x"02200003",x"C83C0008",x"C17DFFFC",x"03DC0020",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0020",x"C05C0014",x"C4240008",x"02200003",x"C83C0008",x"C17DFFFC",x"03DC0020",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0020",x"C05C0014",x"C424000C",x"02200003",x"C83C0008",x"C17DFFFC",x"03DC0020",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0020",x"C05C0014",x"C4240010",x"02200005",x"02600000",x"C17DFFFC",x"00460000",x"03DC0020",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0020",x"02400005",x"02600000",x"C43C0018",x"C17DFFFC",x"00240000",x"00460000",x"03DC0024",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0024",x"02400003",x"C83C0008",x"C43C001C",x"C17DFFFC",x"00240000",x"03DC0028",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0028",x"00420000",x"02200005",x"C17DFFFC",x"03DC0028",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0028",x"02400003",x"C83C0008",x"C43C0020",x"C17DFFFC",x"00240000",x"03DC002C",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC002C",x"C05C0020",x"C4240004",x"02200003",x"C83C0008",x"C17DFFFC",x"03DC002C",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC002C",x"C05C0020",x"C4240008",x"02200003",x"C83C0008",x"C17DFFFC",x"03DC002C",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC002C",x"C05C0020",x"C424000C",x"02200003",x"C83C0008",x"C17DFFFC",x"03DC002C",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC002C",x"C05C0020",x"C4240010",x"02200003",x"C83C0008",x"C17DFFFC",x"03DC002C",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC002C",x"00420000",x"02200005",x"C17DFFFC",x"03DC002C",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC002C",x"02400003",x"C83C0008",x"C43C0024",x"C17DFFFC",x"00240000",x"03DC0030",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0030",x"C05C0024",x"C4240004",x"02200003",x"C83C0008",x"C17DFFFC",x"03DC0030",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0030",x"C05C0024",x"C4240008",x"02200003",x"C83C0008",x"C17DFFFC",x"03DC0030",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0030",x"C05C0024",x"C424000C",x"02200003",x"C83C0008",x"C17DFFFC",x"03DC0030",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0030",x"C05C0024",x"C4240010",x"02200001",x"02600000",x"C17DFFFC",x"00460000",x"03DC0030",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0030",x"02400003",x"C83C0008",x"C43C0028",x"C17DFFFC",x"00240000",x"03DC0034",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0034",x"00420000",x"02200005",x"C17DFFFC",x"03DC0034",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0034",x"02400003",x"C83C0008",x"C43C002C",x"C17DFFFC",x"00240000",x"03DC0038",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0038",x"C05C002C",x"C4240004",x"02200003",x"C83C0008",x"C17DFFFC",x"03DC0038",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0038",x"C05C002C",x"C4240008",x"02200003",x"C83C0008",x"C17DFFFC",x"03DC0038",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0038",x"C05C002C",x"C424000C",x"02200003",x"C83C0008",x"C17DFFFC",x"03DC0038",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0038",x"C05C002C",x"C4240010",x"003A0000",x"03BA0020",x"C442001C",x"C05C0028",x"C4420018",x"C05C0024",x"C4420014",x"C05C0020",x"C4420010",x"C05C001C",x"C442000C",x"C05C0018",x"C4420008",x"C05C0014",x"C4420004",x"C05C0010",x"C4420000",x"C05C0004",x"22640220",x"C09C0000",x"D4286000",x"06240001",x"8620AE08",x"C43C0030",x"C17DFFFC",x"03DC003C",x"037E000C",x"C57DFFFC",x"8200A47C",x"07DC003C",x"C05C0030",x"22640220",x"C09C0000",x"D4286000",x"06440001",x"00280000",x"8200A914",x"00280000",x"C1FDFFFC",x"C1FDFFFC",x"02800005",x"8628AFA0",x"48622000",x"48844000",x"40668000",x"C88000A8",x"40668000",x"C47C0000",x"C45C0004",x"CC5C0008",x"CC3C0010",x"C17DFFFC",x"40206000",x"03DC0020",x"037E000C",x"C57DFFFC",x"8200083C",x"07DC0020",x"CC3C0018",x"C17DFFFC",x"03DC0028",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0028",x"C85C0010",x"48242000",x"C85C0018",x"CC3C0020",x"C17DFFFC",x"40204000",x"03DC0030",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0030",x"C85C0008",x"48242000",x"C85C0018",x"CC3C0028",x"C17DFFFC",x"40204000",x"03DC0038",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0038",x"02200354",x"C05C0004",x"22440220",x"D0224000",x"C05C0000",x"22640220",x"D0626000",x"C0660000",x"C85C0020",x"CC460000",x"C87C0028",x"CC660004",x"CC260008",x"02640028",x"22660220",x"D0626000",x"C0660000",x"44806000",x"CC460000",x"CC260004",x"CC860008",x"02640050",x"22660220",x"D0626000",x"C0660000",x"44A04000",x"CC260000",x"CCA60004",x"CC860008",x"02640001",x"22660220",x"D0626000",x"C0660000",x"44202000",x"CCA60000",x"CC860004",x"CC260008",x"02640029",x"22660220",x"D0626000",x"C0660000",x"CCA60000",x"CC260004",x"CC660008",x"02440051",x"22440220",x"D0224000",x"C0220000",x"CC220000",x"CC420004",x"CC620008",x"C1FDFFFC",x"48244000",x"C840001C",x"40224000",x"C47C0000",x"C45C0004",x"CC9C0030",x"CC5C0038",x"C43C0040",x"CC7C0048",x"C17DFFFC",x"03DC0058",x"037E000C",x"C57DFFFC",x"8200083C",x"07DC0058",x"CC3C0050",x"C17DFFFC",x"03DC0060",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0060",x"C8400068",x"48642000",x"C8800064",x"44668000",x"48662000",x"C8A00060",x"4466A000",x"48662000",x"C8C0005C",x"4066C000",x"48262000",x"C8600058",x"44226000",x"C8FC0048",x"4822E000",x"C9000098",x"CC7C0058",x"CCDC0060",x"CCBC0068",x"CC9C0070",x"CC5C0078",x"CD1C0080",x"CC3C0088",x"8E30B07C",x"45230000",x"C17DFFFC",x"40212000",x"03DC0098",x"037E000C",x"C57DFFFC",x"82000EC4",x"07DC0098",x"8200B0E8",x"8E02B0CC",x"C9200090",x"8F22B0AC",x"41230000",x"C17DFFFC",x"40212000",x"03DC0098",x"037E000C",x"C57DFFFC",x"82000EC4",x"07DC0098",x"8200B0C8",x"02200001",x"C17DFFFC",x"03DC0098",x"037E000C",x"C57DFFFC",x"8200084C",x"07DC0098",x"8200B0E8",x"0220FFFF",x"C17DFFFC",x"03DC0098",x"037E000C",x"C57DFFFC",x"8200084C",x"07DC0098",x"C85C0080",x"C87C0088",x"CC3C0090",x"8E64B11C",x"44664000",x"C17DFFFC",x"40206000",x"03DC00A0",x"037E000C",x"C57DFFFC",x"82001270",x"07DC00A0",x"8200B190",x"8E06B170",x"C8800090",x"8E86B14C",x"40664000",x"C17DFFFC",x"40206000",x"03DC00A0",x"037E000C",x"C57DFFFC",x"82001270",x"07DC00A0",x"8200B16C",x"02200001",x"C17DFFFC",x"40206000",x"03DC00A0",x"037E000C",x"C57DFFFC",x"82000B88",x"07DC00A0",x"8200B190",x"0220FFFF",x"C17DFFFC",x"40206000",x"03DC00A0",x"037E000C",x"C57DFFFC",x"82000B88",x"07DC00A0",x"C17DFFFC",x"03DC00A0",x"037E000C",x"C57DFFFC",x"82000844",x"07DC00A0",x"C85C0090",x"48242000",x"C85C0050",x"48224000",x"C03C0040",x"02220001",x"48422000",x"C87C0038",x"40446000",x"CC3C0098",x"C43C00A0",x"C17DFFFC",x"40204000",x"03DC00AC",x"037E000C",x"C57DFFFC",x"8200083C",x"07DC00AC",x"CC3C00A8",x"C17DFFFC",x"03DC00B8",x"037E000C",x"C57DFFFC",x"82000844",x"07DC00B8",x"C85C0078",x"48442000",x"C87C0070",x"44446000",x"48442000",x"C87C0068",x"44446000",x"48442000",x"C87C0060",x"40446000",x"48242000",x"C85C0058",x"44224000",x"C85C0030",x"48224000",x"C87C0080",x"CC3C00B0",x"8E26B278",x"44826000",x"C17DFFFC",x"40208000",x"03DC00C0",x"037E000C",x"C57DFFFC",x"82000EC4",x"07DC00C0",x"8200B2E4",x"8E02B2C8",x"C8800090",x"8E82B2A8",x"40826000",x"C17DFFFC",x"40208000",x"03DC00C0",x"037E000C",x"C57DFFFC",x"82000EC4",x"07DC00C0",x"8200B2C4",x"02200001",x"C17DFFFC",x"03DC00C0",x"037E000C",x"C57DFFFC",x"8200084C",x"07DC00C0",x"8200B2E4",x"0220FFFF",x"C17DFFFC",x"03DC00C0",x"037E000C",x"C57DFFFC",x"8200084C",x"07DC00C0",x"C85C0080",x"C87C00B0",x"CC3C00B8",x"8E64B318",x"44464000",x"C17DFFFC",x"40204000",x"03DC00C8",x"037E000C",x"C57DFFFC",x"82001270",x"07DC00C8",x"8200B38C",x"8E06B36C",x"C8800090",x"8E86B348",x"40464000",x"C17DFFFC",x"40204000",x"03DC00C8",x"037E000C",x"C57DFFFC",x"82001270",x"07DC00C8",x"8200B368",x"02200001",x"C17DFFFC",x"40206000",x"03DC00C8",x"037E000C",x"C57DFFFC",x"82000B88",x"07DC00C8",x"8200B38C",x"0220FFFF",x"C17DFFFC",x"40206000",x"03DC00C8",x"037E000C",x"C57DFFFC",x"82000B88",x"07DC00C8",x"C17DFFFC",x"03DC00C8",x"037E000C",x"C57DFFFC",x"82000844",x"07DC00C8",x"C85C00B8",x"48242000",x"C85C00A8",x"48424000",x"C83C0098",x"C87C0048",x"C89C0030",x"C03C00A0",x"C05C0004",x"C07C0000",x"8200AE14",x"8620B570",x"58420000",x"C8600010",x"48446000",x"C880000C",x"44A48000",x"02800000",x"40C00000",x"CC9C0000",x"CC7C0008",x"C43C0010",x"CC3C0018",x"CCDC0020",x"C45C0028",x"C47C002C",x"CC5C0030",x"C17DFFFC",x"00280000",x"40802000",x"4060A000",x"4040C000",x"4020C000",x"03DC0040",x"037E000C",x"C57DFFFC",x"8200AE14",x"07DC0040",x"C820001C",x"C85C0030",x"40642000",x"02200000",x"C05C002C",x"02640002",x"C85C0020",x"C89C0018",x"C09C0028",x"CC3C0038",x"C17DFFFC",x"00480000",x"40204000",x"03DC0048",x"037E000C",x"C57DFFFC",x"8200AE14",x"07DC0048",x"C03C0010",x"06220001",x"C05C0028",x"02440001",x"02600005",x"8646B4A4",x"06440005",x"8200B4A4",x"8620B56C",x"58220000",x"C85C0008",x"48224000",x"C85C0000",x"44624000",x"02600000",x"C85C0020",x"C89C0018",x"C09C002C",x"C43C0040",x"C45C0044",x"CC3C0048",x"C17DFFFC",x"00260000",x"00680000",x"40204000",x"03DC0058",x"037E000C",x"C57DFFFC",x"8200AE14",x"07DC0058",x"C83C0038",x"C85C0048",x"40642000",x"02200000",x"C05C002C",x"02640002",x"C83C0020",x"C89C0018",x"C09C0044",x"C17DFFFC",x"00480000",x"40402000",x"03DC0058",x"037E000C",x"C57DFFFC",x"8200AE14",x"07DC0058",x"C03C0040",x"06220001",x"C05C0044",x"02440001",x"02600005",x"8646B560",x"06440005",x"8200B560",x"C83C0018",x"C07C002C",x"8200B3D0",x"C1FDFFFC",x"C1FDFFFC",x"8620B6F8",x"58220000",x"C8400010",x"48224000",x"C860000C",x"44826000",x"C8200008",x"02800000",x"40A00000",x"CC5C0000",x"C43C0008",x"CC9C0010",x"CC7C0018",x"CCBC0020",x"C45C0028",x"C47C002C",x"C17DFFFC",x"00280000",x"40602000",x"4040A000",x"4020A000",x"03DC0038",x"037E000C",x"C57DFFFC",x"8200AE14",x"07DC0038",x"02200000",x"C05C002C",x"02640002",x"C83C0020",x"C87C0018",x"C89C0010",x"C09C0028",x"C17DFFFC",x"00480000",x"40402000",x"03DC0038",x"037E000C",x"C57DFFFC",x"8200AE14",x"07DC0038",x"02200003",x"C05C0028",x"02640001",x"02800005",x"8668B634",x"06660005",x"8200B634",x"C83C0010",x"C09C002C",x"C17DFFFC",x"00460000",x"00680000",x"03DC0038",x"037E000C",x"C57DFFFC",x"8200B3D0",x"07DC0038",x"C03C0008",x"06220001",x"C05C0028",x"02440002",x"02600005",x"8646B67C",x"06440005",x"8200B67C",x"C07C002C",x"02660004",x"8620B6F4",x"58220000",x"C85C0000",x"48224000",x"C85C0018",x"44224000",x"02800004",x"C47C0030",x"C45C0034",x"C43C0038",x"C17DFFFC",x"00280000",x"03DC0044",x"037E000C",x"C57DFFFC",x"8200B3D0",x"07DC0044",x"C03C0038",x"06220001",x"C05C0034",x"02440002",x"02600005",x"8646B6E8",x"06440005",x"8200B6E8",x"C07C0030",x"02660004",x"8200B574",x"C1FDFFFC",x"C1FDFFFC",x"8640B928",x"02600003",x"40200000",x"CC3C0000",x"C43C0008",x"C45C000C",x"C17DFFFC",x"00260000",x"03DC0018",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0018",x"00420000",x"022000C4",x"C0620000",x"C43C0010",x"C45C0014",x"C17DFFFC",x"00260000",x"03DC0020",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0020",x"005A0000",x"03BA0008",x"C4240004",x"C03C0014",x"C4240000",x"00240000",x"C05C000C",x"22640220",x"C09C0008",x"D4286000",x"06240001",x"8620B924",x"02400003",x"C83C0000",x"C43C0018",x"C17DFFFC",x"00240000",x"03DC0024",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0024",x"00420000",x"C03C0010",x"C0620000",x"C45C001C",x"C17DFFFC",x"00260000",x"03DC0028",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0028",x"005A0000",x"03BA0008",x"C4240004",x"C03C001C",x"C4240000",x"00240000",x"C05C0018",x"22640220",x"C09C0008",x"D4286000",x"06240001",x"8620B920",x"02400003",x"C83C0000",x"C43C0020",x"C17DFFFC",x"00240000",x"03DC002C",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC002C",x"00420000",x"C03C0010",x"C0620000",x"C45C0024",x"C17DFFFC",x"00260000",x"03DC0030",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0030",x"005A0000",x"03BA0008",x"C4240004",x"C03C0024",x"C4240000",x"00240000",x"C05C0020",x"22640220",x"C09C0008",x"D4286000",x"06240001",x"8620B91C",x"02400003",x"C83C0000",x"C43C0028",x"C17DFFFC",x"00240000",x"03DC0034",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0034",x"00420000",x"C03C0010",x"C0220000",x"C45C002C",x"C17DFFFC",x"03DC0038",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0038",x"005A0000",x"03BA0008",x"C4240004",x"C03C002C",x"C4240000",x"00240000",x"C05C0028",x"22640220",x"C09C0008",x"D4286000",x"06440001",x"00280000",x"8200B6FC",x"C1FDFFFC",x"C1FDFFFC",x"C1FDFFFC",x"C1FDFFFC",x"8620BD0C",x"02400354",x"02600078",x"02800003",x"40200000",x"CC3C0000",x"C45C0008",x"C43C000C",x"C47C0010",x"C17DFFFC",x"00280000",x"03DC001C",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC001C",x"00420000",x"022000C4",x"C0620000",x"C43C0014",x"C45C0018",x"C17DFFFC",x"00260000",x"03DC0024",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0024",x"005A0000",x"03BA0008",x"C4240004",x"C03C0018",x"C4240000",x"C03C0010",x"C17DFFFC",x"03DC0024",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0024",x"C05C000C",x"22640220",x"C09C0008",x"D4286000",x"02600003",x"C83C0000",x"C43C001C",x"C17DFFFC",x"00260000",x"03DC0028",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0028",x"00420000",x"C03C0014",x"C0620000",x"C45C0020",x"C17DFFFC",x"00260000",x"03DC002C",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC002C",x"005A0000",x"03BA0008",x"C4240004",x"C03C0020",x"C4240000",x"00240000",x"C05C001C",x"C42401D8",x"02200003",x"C83C0000",x"C17DFFFC",x"03DC002C",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC002C",x"00420000",x"C03C0014",x"C0620000",x"C45C0024",x"C17DFFFC",x"00260000",x"03DC0030",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0030",x"005A0000",x"03BA0008",x"C4240004",x"C03C0024",x"C4240000",x"00240000",x"C05C001C",x"C42401D4",x"02200003",x"C83C0000",x"C17DFFFC",x"03DC0030",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0030",x"00420000",x"C03C0014",x"C0620000",x"C45C0028",x"C17DFFFC",x"00260000",x"03DC0034",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0034",x"005A0000",x"03BA0008",x"C4240004",x"C03C0028",x"C4240000",x"00240000",x"C05C001C",x"C42401D0",x"02200073",x"C17DFFFC",x"01240000",x"00420000",x"00320000",x"03DC0034",x"037E000C",x"C57DFFFC",x"8200B6FC",x"07DC0034",x"C03C000C",x"06220001",x"8620BD08",x"02400078",x"02600003",x"C83C0000",x"C43C002C",x"C45C0030",x"C17DFFFC",x"00260000",x"03DC003C",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC003C",x"00420000",x"C03C0014",x"C0620000",x"C45C0034",x"C17DFFFC",x"00260000",x"03DC0040",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0040",x"005A0000",x"03BA0008",x"C4240004",x"C03C0034",x"C4240000",x"C03C0030",x"C17DFFFC",x"03DC0040",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0040",x"C05C002C",x"22640220",x"C09C0008",x"D4286000",x"02600003",x"C83C0000",x"C43C0038",x"C17DFFFC",x"00260000",x"03DC0044",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0044",x"00420000",x"C03C0014",x"C0620000",x"C45C003C",x"C17DFFFC",x"00260000",x"03DC0048",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0048",x"005A0000",x"03BA0008",x"C4240004",x"C03C003C",x"C4240000",x"00240000",x"C05C0038",x"C42401D8",x"02200003",x"C83C0000",x"C17DFFFC",x"03DC0048",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0048",x"00420000",x"C03C0014",x"C0220000",x"C45C0040",x"C17DFFFC",x"03DC004C",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC004C",x"005A0000",x"03BA0008",x"C4240004",x"C03C0040",x"C4240000",x"00240000",x"C05C0038",x"C42401D4",x"02200074",x"C17DFFFC",x"01240000",x"00420000",x"00320000",x"03DC004C",x"037E000C",x"C57DFFFC",x"8200B6FC",x"07DC004C",x"C03C002C",x"06220001",x"8200B92C",x"C1FDFFFC",x"C1FDFFFC",x"8640C710",x"22640220",x"D0626000",x"028000C4",x"C0A80000",x"06AA0001",x"C49C0000",x"C43C0004",x"C45C0008",x"86A0BF18",x"02C000C8",x"22EA0220",x"D0ECE000",x"C1060004",x"C1260000",x"C14E0004",x"02800001",x"C47C000C",x"C4DC0010",x"8348BDE0",x"02800002",x"8348BDA4",x"C51C0014",x"C4BC0018",x"C17DFFFC",x"004E0000",x"00320000",x"03DC0024",x"037E000C",x"C57DFFFC",x"8200400C",x"07DC0024",x"C05C0018",x"22640220",x"C09C0014",x"D4286000",x"8200BDDC",x"C51C0014",x"C4BC0018",x"C17DFFFC",x"004E0000",x"00320000",x"03DC0024",x"037E000C",x"C57DFFFC",x"82003E98",x"07DC0024",x"C05C0018",x"22640220",x"C09C0014",x"D4286000",x"8200BE18",x"C51C0014",x"C4BC0018",x"C17DFFFC",x"004E0000",x"00320000",x"03DC0024",x"037E000C",x"C57DFFFC",x"82003CC4",x"07DC0024",x"C05C0018",x"22640220",x"C09C0014",x"D4286000",x"06240001",x"8620BF14",x"22420220",x"C07C0010",x"D0464000",x"C07C000C",x"C0860004",x"C0A60000",x"C0C40004",x"02E00001",x"82CEBEBC",x"02E00002",x"82CEBE84",x"C49C001C",x"C43C0020",x"C17DFFFC",x"002A0000",x"03DC002C",x"037E000C",x"C57DFFFC",x"8200400C",x"07DC002C",x"C05C0020",x"22640220",x"C09C001C",x"D4286000",x"8200BEB8",x"C49C001C",x"C43C0020",x"C17DFFFC",x"002A0000",x"03DC002C",x"037E000C",x"C57DFFFC",x"82003E98",x"07DC002C",x"C05C0020",x"22640220",x"C09C001C",x"D4286000",x"8200BEF0",x"C49C001C",x"C43C0020",x"C17DFFFC",x"002A0000",x"03DC002C",x"037E000C",x"C57DFFFC",x"82003CC4",x"07DC002C",x"C05C0020",x"22640220",x"C09C001C",x"D4286000",x"06440001",x"C03C000C",x"C17DFFFC",x"03DC002C",x"037E000C",x"C57DFFFC",x"820042A4",x"07DC002C",x"8200BF14",x"8200BF18",x"C03C0008",x"06220001",x"8620C70C",x"22420220",x"C07C0004",x"D0464000",x"C09C0000",x"C0A80000",x"06AA0001",x"C43C0024",x"86A0C200",x"02C000C8",x"22EA0220",x"D0ECE000",x"C1040004",x"C1240000",x"C14E0004",x"02800001",x"C45C0028",x"C4DC002C",x"8348BFEC",x"02800002",x"8348BFB0",x"C51C0030",x"C4BC0034",x"C17DFFFC",x"004E0000",x"00320000",x"03DC0040",x"037E000C",x"C57DFFFC",x"8200400C",x"07DC0040",x"C05C0034",x"22640220",x"C09C0030",x"D4286000",x"8200BFE8",x"C51C0030",x"C4BC0034",x"C17DFFFC",x"004E0000",x"00320000",x"03DC0040",x"037E000C",x"C57DFFFC",x"82003E98",x"07DC0040",x"C05C0034",x"22640220",x"C09C0030",x"D4286000",x"8200C024",x"C51C0030",x"C4BC0034",x"C17DFFFC",x"004E0000",x"00320000",x"03DC0040",x"037E000C",x"C57DFFFC",x"82003CC4",x"07DC0040",x"C05C0034",x"22640220",x"C09C0030",x"D4286000",x"06240001",x"8620C1FC",x"22420220",x"C07C002C",x"D0464000",x"C09C0028",x"C0A80004",x"C0C80000",x"C0E40004",x"03000001",x"82F0C0C8",x"03000002",x"82F0C090",x"C4BC0038",x"C43C003C",x"C17DFFFC",x"002C0000",x"03DC0048",x"037E000C",x"C57DFFFC",x"8200400C",x"07DC0048",x"C05C003C",x"22640220",x"C09C0038",x"D4286000",x"8200C0C4",x"C4BC0038",x"C43C003C",x"C17DFFFC",x"002C0000",x"03DC0048",x"037E000C",x"C57DFFFC",x"82003E98",x"07DC0048",x"C05C003C",x"22640220",x"C09C0038",x"D4286000",x"8200C0FC",x"C4BC0038",x"C43C003C",x"C17DFFFC",x"002C0000",x"03DC0048",x"037E000C",x"C57DFFFC",x"82003CC4",x"07DC0048",x"C05C003C",x"22640220",x"C09C0038",x"D4286000",x"06240001",x"8620C1F8",x"22420220",x"C07C002C",x"D0464000",x"C07C0028",x"C0860004",x"C0A60000",x"C0C40004",x"02E00001",x"82CEC1A0",x"02E00002",x"82CEC168",x"C49C0040",x"C43C0044",x"C17DFFFC",x"002A0000",x"03DC0050",x"037E000C",x"C57DFFFC",x"8200400C",x"07DC0050",x"C05C0044",x"22640220",x"C09C0040",x"D4286000",x"8200C19C",x"C49C0040",x"C43C0044",x"C17DFFFC",x"002A0000",x"03DC0050",x"037E000C",x"C57DFFFC",x"82003E98",x"07DC0050",x"C05C0044",x"22640220",x"C09C0040",x"D4286000",x"8200C1D4",x"C49C0040",x"C43C0044",x"C17DFFFC",x"002A0000",x"03DC0050",x"037E000C",x"C57DFFFC",x"82003CC4",x"07DC0050",x"C05C0044",x"22640220",x"C09C0040",x"D4286000",x"06440001",x"C03C0028",x"C17DFFFC",x"03DC0050",x"037E000C",x"C57DFFFC",x"820042A4",x"07DC0050",x"8200C1F8",x"8200C1FC",x"8200C200",x"C03C0024",x"06220001",x"8620C708",x"22420220",x"C07C0004",x"D0464000",x"C09C0000",x"C0A80000",x"06AA0001",x"C43C0048",x"86A0C40C",x"02C000C8",x"22EA0220",x"D0ECE000",x"C1040004",x"C1240000",x"C14E0004",x"02800001",x"C45C004C",x"C4DC0050",x"8348C2D4",x"02800002",x"8348C298",x"C51C0054",x"C4BC0058",x"C17DFFFC",x"004E0000",x"00320000",x"03DC0064",x"037E000C",x"C57DFFFC",x"8200400C",x"07DC0064",x"C05C0058",x"22640220",x"C09C0054",x"D4286000",x"8200C2D0",x"C51C0054",x"C4BC0058",x"C17DFFFC",x"004E0000",x"00320000",x"03DC0064",x"037E000C",x"C57DFFFC",x"82003E98",x"07DC0064",x"C05C0058",x"22640220",x"C09C0054",x"D4286000",x"8200C30C",x"C51C0054",x"C4BC0058",x"C17DFFFC",x"004E0000",x"00320000",x"03DC0064",x"037E000C",x"C57DFFFC",x"82003CC4",x"07DC0064",x"C05C0058",x"22640220",x"C09C0054",x"D4286000",x"06240001",x"8620C408",x"22420220",x"C07C0050",x"D0464000",x"C07C004C",x"C0860004",x"C0A60000",x"C0C40004",x"02E00001",x"82CEC3B0",x"02E00002",x"82CEC378",x"C49C005C",x"C43C0060",x"C17DFFFC",x"002A0000",x"03DC006C",x"037E000C",x"C57DFFFC",x"8200400C",x"07DC006C",x"C05C0060",x"22640220",x"C09C005C",x"D4286000",x"8200C3AC",x"C49C005C",x"C43C0060",x"C17DFFFC",x"002A0000",x"03DC006C",x"037E000C",x"C57DFFFC",x"82003E98",x"07DC006C",x"C05C0060",x"22640220",x"C09C005C",x"D4286000",x"8200C3E4",x"C49C005C",x"C43C0060",x"C17DFFFC",x"002A0000",x"03DC006C",x"037E000C",x"C57DFFFC",x"82003CC4",x"07DC006C",x"C05C0060",x"22640220",x"C09C005C",x"D4286000",x"06440001",x"C03C004C",x"C17DFFFC",x"03DC006C",x"037E000C",x"C57DFFFC",x"820042A4",x"07DC006C",x"8200C408",x"8200C40C",x"C03C0048",x"06220001",x"8620C704",x"22420220",x"C07C0004",x"D0464000",x"C09C0000",x"C0880000",x"06880001",x"C43C0064",x"8680C6F4",x"02A000C8",x"22C80220",x"D0CAC000",x"C0E40004",x"C1040000",x"C12C0004",x"03400001",x"C45C0068",x"C4BC006C",x"8334C4E0",x"03400002",x"8334C4A4",x"C4FC0070",x"C49C0074",x"C17DFFFC",x"004C0000",x"00300000",x"03DC0080",x"037E000C",x"C57DFFFC",x"8200400C",x"07DC0080",x"C05C0074",x"22640220",x"C09C0070",x"D4286000",x"8200C4DC",x"C4FC0070",x"C49C0074",x"C17DFFFC",x"004C0000",x"00300000",x"03DC0080",x"037E000C",x"C57DFFFC",x"82003E98",x"07DC0080",x"C05C0074",x"22640220",x"C09C0070",x"D4286000",x"8200C518",x"C4FC0070",x"C49C0074",x"C17DFFFC",x"004C0000",x"00300000",x"03DC0080",x"037E000C",x"C57DFFFC",x"82003CC4",x"07DC0080",x"C05C0074",x"22640220",x"C09C0070",x"D4286000",x"06240001",x"8620C6F0",x"22420220",x"C07C006C",x"D0464000",x"C09C0068",x"C0A80004",x"C0C80000",x"C0E40004",x"03000001",x"82F0C5BC",x"03000002",x"82F0C584",x"C4BC0078",x"C43C007C",x"C17DFFFC",x"002C0000",x"03DC0088",x"037E000C",x"C57DFFFC",x"8200400C",x"07DC0088",x"C05C007C",x"22640220",x"C09C0078",x"D4286000",x"8200C5B8",x"C4BC0078",x"C43C007C",x"C17DFFFC",x"002C0000",x"03DC0088",x"037E000C",x"C57DFFFC",x"82003E98",x"07DC0088",x"C05C007C",x"22640220",x"C09C0078",x"D4286000",x"8200C5F0",x"C4BC0078",x"C43C007C",x"C17DFFFC",x"002C0000",x"03DC0088",x"037E000C",x"C57DFFFC",x"82003CC4",x"07DC0088",x"C05C007C",x"22640220",x"C09C0078",x"D4286000",x"06240001",x"8620C6EC",x"22420220",x"C07C006C",x"D0464000",x"C07C0068",x"C0860004",x"C0A60000",x"C0C40004",x"02E00001",x"82CEC694",x"02E00002",x"82CEC65C",x"C49C0080",x"C43C0084",x"C17DFFFC",x"002A0000",x"03DC0090",x"037E000C",x"C57DFFFC",x"8200400C",x"07DC0090",x"C05C0084",x"22640220",x"C09C0080",x"D4286000",x"8200C690",x"C49C0080",x"C43C0084",x"C17DFFFC",x"002A0000",x"03DC0090",x"037E000C",x"C57DFFFC",x"82003E98",x"07DC0090",x"C05C0084",x"22640220",x"C09C0080",x"D4286000",x"8200C6C8",x"C49C0080",x"C43C0084",x"C17DFFFC",x"002A0000",x"03DC0090",x"037E000C",x"C57DFFFC",x"82003CC4",x"07DC0090",x"C05C0084",x"22640220",x"C09C0080",x"D4286000",x"06440001",x"C03C0068",x"C17DFFFC",x"03DC0090",x"037E000C",x"C57DFFFC",x"820042A4",x"07DC0090",x"8200C6EC",x"8200C6F0",x"8200C6F4",x"C03C0064",x"06420001",x"C03C0004",x"8200BD10",x"C1FDFFFC",x"C1FDFFFC",x"C1FDFFFC",x"C1FDFFFC",x"8620D760",x"02400354",x"22620220",x"D0646000",x"C08601DC",x"02A000C4",x"C0CA0000",x"06CC0001",x"C45C0000",x"C43C0004",x"C4BC0008",x"C47C000C",x"86C0CA04",x"02E000C8",x"230C0220",x"D10F0000",x"C1280004",x"C1480000",x"C0500004",x"02200001",x"C49C0010",x"C4FC0014",x"8242C7F0",x"02200002",x"8242C7B4",x"C53C0018",x"C4DC001C",x"C17DFFFC",x"00500000",x"00340000",x"03DC0028",x"037E000C",x"C57DFFFC",x"8200400C",x"07DC0028",x"C05C001C",x"22640220",x"C09C0018",x"D4286000",x"8200C7EC",x"C53C0018",x"C4DC001C",x"C17DFFFC",x"00500000",x"00340000",x"03DC0028",x"037E000C",x"C57DFFFC",x"82003E98",x"07DC0028",x"C05C001C",x"22640220",x"C09C0018",x"D4286000",x"8200C828",x"C53C0018",x"C4DC001C",x"C17DFFFC",x"00500000",x"00340000",x"03DC0028",x"037E000C",x"C57DFFFC",x"82003CC4",x"07DC0028",x"C05C001C",x"22640220",x"C09C0018",x"D4286000",x"06240001",x"8620CA00",x"22420220",x"C07C0014",x"D0464000",x"C09C0010",x"C0A80004",x"C0C80000",x"C0E40004",x"03000001",x"82F0C8CC",x"03000002",x"82F0C894",x"C4BC0020",x"C43C0024",x"C17DFFFC",x"002C0000",x"03DC0030",x"037E000C",x"C57DFFFC",x"8200400C",x"07DC0030",x"C05C0024",x"22640220",x"C09C0020",x"D4286000",x"8200C8C8",x"C4BC0020",x"C43C0024",x"C17DFFFC",x"002C0000",x"03DC0030",x"037E000C",x"C57DFFFC",x"82003E98",x"07DC0030",x"C05C0024",x"22640220",x"C09C0020",x"D4286000",x"8200C900",x"C4BC0020",x"C43C0024",x"C17DFFFC",x"002C0000",x"03DC0030",x"037E000C",x"C57DFFFC",x"82003CC4",x"07DC0030",x"C05C0024",x"22640220",x"C09C0020",x"D4286000",x"06240001",x"8620C9FC",x"22420220",x"C07C0014",x"D0464000",x"C07C0010",x"C0860004",x"C0A60000",x"C0C40004",x"02E00001",x"82CEC9A4",x"02E00002",x"82CEC96C",x"C49C0028",x"C43C002C",x"C17DFFFC",x"002A0000",x"03DC0038",x"037E000C",x"C57DFFFC",x"8200400C",x"07DC0038",x"C05C002C",x"22640220",x"C09C0028",x"D4286000",x"8200C9A0",x"C49C0028",x"C43C002C",x"C17DFFFC",x"002A0000",x"03DC0038",x"037E000C",x"C57DFFFC",x"82003E98",x"07DC0038",x"C05C002C",x"22640220",x"C09C0028",x"D4286000",x"8200C9D8",x"C49C0028",x"C43C002C",x"C17DFFFC",x"002A0000",x"03DC0038",x"037E000C",x"C57DFFFC",x"82003CC4",x"07DC0038",x"C05C002C",x"22640220",x"C09C0028",x"D4286000",x"06440001",x"C03C0010",x"C17DFFFC",x"03DC0038",x"037E000C",x"C57DFFFC",x"820042A4",x"07DC0038",x"8200C9FC",x"8200CA00",x"8200CA04",x"C03C000C",x"C04201D8",x"C07C0008",x"C0860000",x"06880001",x"8680CBFC",x"02A000C8",x"22C80220",x"D0CAC000",x"C0E40004",x"C1040000",x"C12C0004",x"03400001",x"C45C0030",x"C4BC0034",x"8334CAC4",x"03400002",x"8334CA88",x"C4FC0038",x"C49C003C",x"C17DFFFC",x"004C0000",x"00300000",x"03DC0048",x"037E000C",x"C57DFFFC",x"8200400C",x"07DC0048",x"C05C003C",x"22640220",x"C09C0038",x"D4286000",x"8200CAC0",x"C4FC0038",x"C49C003C",x"C17DFFFC",x"004C0000",x"00300000",x"03DC0048",x"037E000C",x"C57DFFFC",x"82003E98",x"07DC0048",x"C05C003C",x"22640220",x"C09C0038",x"D4286000",x"8200CAFC",x"C4FC0038",x"C49C003C",x"C17DFFFC",x"004C0000",x"00300000",x"03DC0048",x"037E000C",x"C57DFFFC",x"82003CC4",x"07DC0048",x"C05C003C",x"22640220",x"C09C0038",x"D4286000",x"06240001",x"8620CBF8",x"22420220",x"C07C0034",x"D0464000",x"C07C0030",x"C0860004",x"C0A60000",x"C0C40004",x"02E00001",x"82CECBA0",x"02E00002",x"82CECB68",x"C49C0040",x"C43C0044",x"C17DFFFC",x"002A0000",x"03DC0050",x"037E000C",x"C57DFFFC",x"8200400C",x"07DC0050",x"C05C0044",x"22640220",x"C09C0040",x"D4286000",x"8200CB9C",x"C49C0040",x"C43C0044",x"C17DFFFC",x"002A0000",x"03DC0050",x"037E000C",x"C57DFFFC",x"82003E98",x"07DC0050",x"C05C0044",x"22640220",x"C09C0040",x"D4286000",x"8200CBD4",x"C49C0040",x"C43C0044",x"C17DFFFC",x"002A0000",x"03DC0050",x"037E000C",x"C57DFFFC",x"82003CC4",x"07DC0050",x"C05C0044",x"22640220",x"C09C0040",x"D4286000",x"06440001",x"C03C0030",x"C17DFFFC",x"03DC0050",x"037E000C",x"C57DFFFC",x"820042A4",x"07DC0050",x"8200CBF8",x"8200CBFC",x"C03C000C",x"C04201D4",x"C07C0008",x"C0860000",x"06880001",x"8680CED0",x"02A000C8",x"22C80220",x"D0CAC000",x"C0E40004",x"C1040000",x"C12C0004",x"03400001",x"C45C0048",x"C4BC004C",x"8334CCBC",x"03400002",x"8334CC80",x"C4FC0050",x"C49C0054",x"C17DFFFC",x"004C0000",x"00300000",x"03DC0060",x"037E000C",x"C57DFFFC",x"8200400C",x"07DC0060",x"C05C0054",x"22640220",x"C09C0050",x"D4286000",x"8200CCB8",x"C4FC0050",x"C49C0054",x"C17DFFFC",x"004C0000",x"00300000",x"03DC0060",x"037E000C",x"C57DFFFC",x"82003E98",x"07DC0060",x"C05C0054",x"22640220",x"C09C0050",x"D4286000",x"8200CCF4",x"C4FC0050",x"C49C0054",x"C17DFFFC",x"004C0000",x"00300000",x"03DC0060",x"037E000C",x"C57DFFFC",x"82003CC4",x"07DC0060",x"C05C0054",x"22640220",x"C09C0050",x"D4286000",x"06240001",x"8620CECC",x"22420220",x"C07C004C",x"D0464000",x"C09C0048",x"C0A80004",x"C0C80000",x"C0E40004",x"03000001",x"82F0CD98",x"03000002",x"82F0CD60",x"C4BC0058",x"C43C005C",x"C17DFFFC",x"002C0000",x"03DC0068",x"037E000C",x"C57DFFFC",x"8200400C",x"07DC0068",x"C05C005C",x"22640220",x"C09C0058",x"D4286000",x"8200CD94",x"C4BC0058",x"C43C005C",x"C17DFFFC",x"002C0000",x"03DC0068",x"037E000C",x"C57DFFFC",x"82003E98",x"07DC0068",x"C05C005C",x"22640220",x"C09C0058",x"D4286000",x"8200CDCC",x"C4BC0058",x"C43C005C",x"C17DFFFC",x"002C0000",x"03DC0068",x"037E000C",x"C57DFFFC",x"82003CC4",x"07DC0068",x"C05C005C",x"22640220",x"C09C0058",x"D4286000",x"06240001",x"8620CEC8",x"22420220",x"C07C004C",x"D0464000",x"C07C0048",x"C0860004",x"C0A60000",x"C0C40004",x"02E00001",x"82CECE70",x"02E00002",x"82CECE38",x"C49C0060",x"C43C0064",x"C17DFFFC",x"002A0000",x"03DC0070",x"037E000C",x"C57DFFFC",x"8200400C",x"07DC0070",x"C05C0064",x"22640220",x"C09C0060",x"D4286000",x"8200CE6C",x"C49C0060",x"C43C0064",x"C17DFFFC",x"002A0000",x"03DC0070",x"037E000C",x"C57DFFFC",x"82003E98",x"07DC0070",x"C05C0064",x"22640220",x"C09C0060",x"D4286000",x"8200CEA4",x"C49C0060",x"C43C0064",x"C17DFFFC",x"002A0000",x"03DC0070",x"037E000C",x"C57DFFFC",x"82003CC4",x"07DC0070",x"C05C0064",x"22640220",x"C09C0060",x"D4286000",x"06440001",x"C03C0048",x"C17DFFFC",x"03DC0070",x"037E000C",x"C57DFFFC",x"820042A4",x"07DC0070",x"8200CEC8",x"8200CECC",x"8200CED0",x"02400074",x"C03C000C",x"C17DFFFC",x"03DC0070",x"037E000C",x"C57DFFFC",x"8200BD10",x"07DC0070",x"C03C0004",x"06220001",x"8620D75C",x"22420220",x"C07C0000",x"D0464000",x"C08401DC",x"C0BC0008",x"C0CA0000",x"06CC0001",x"C43C0068",x"C45C006C",x"86C0D104",x"02E000C8",x"230C0220",x"D10F0000",x"C1280004",x"C1480000",x"C0700004",x"02200001",x"C49C0070",x"C4FC0074",x"8262CFCC",x"02200002",x"8262CF90",x"C53C0078",x"C4DC007C",x"C17DFFFC",x"00500000",x"00340000",x"03DC0088",x"037E000C",x"C57DFFFC",x"8200400C",x"07DC0088",x"C05C007C",x"22640220",x"C09C0078",x"D4286000",x"8200CFC8",x"C53C0078",x"C4DC007C",x"C17DFFFC",x"00500000",x"00340000",x"03DC0088",x"037E000C",x"C57DFFFC",x"82003E98",x"07DC0088",x"C05C007C",x"22640220",x"C09C0078",x"D4286000",x"8200D004",x"C53C0078",x"C4DC007C",x"C17DFFFC",x"00500000",x"00340000",x"03DC0088",x"037E000C",x"C57DFFFC",x"82003CC4",x"07DC0088",x"C05C007C",x"22640220",x"C09C0078",x"D4286000",x"06240001",x"8620D100",x"22420220",x"C07C0074",x"D0464000",x"C07C0070",x"C0860004",x"C0A60000",x"C0C40004",x"02E00001",x"82CED0A8",x"02E00002",x"82CED070",x"C49C0080",x"C43C0084",x"C17DFFFC",x"002A0000",x"03DC0090",x"037E000C",x"C57DFFFC",x"8200400C",x"07DC0090",x"C05C0084",x"22640220",x"C09C0080",x"D4286000",x"8200D0A4",x"C49C0080",x"C43C0084",x"C17DFFFC",x"002A0000",x"03DC0090",x"037E000C",x"C57DFFFC",x"82003E98",x"07DC0090",x"C05C0084",x"22640220",x"C09C0080",x"D4286000",x"8200D0DC",x"C49C0080",x"C43C0084",x"C17DFFFC",x"002A0000",x"03DC0090",x"037E000C",x"C57DFFFC",x"82003CC4",x"07DC0090",x"C05C0084",x"22640220",x"C09C0080",x"D4286000",x"06440001",x"C03C0070",x"C17DFFFC",x"03DC0090",x"037E000C",x"C57DFFFC",x"820042A4",x"07DC0090",x"8200D100",x"8200D104",x"C03C006C",x"C04201D8",x"C07C0008",x"C0860000",x"06880001",x"8680D3D8",x"02A000C8",x"22C80220",x"D0CAC000",x"C0E40004",x"C1040000",x"C12C0004",x"03400001",x"C45C0088",x"C4BC008C",x"8334D1C4",x"03400002",x"8334D188",x"C4FC0090",x"C49C0094",x"C17DFFFC",x"004C0000",x"00300000",x"03DC00A0",x"037E000C",x"C57DFFFC",x"8200400C",x"07DC00A0",x"C05C0094",x"22640220",x"C09C0090",x"D4286000",x"8200D1C0",x"C4FC0090",x"C49C0094",x"C17DFFFC",x"004C0000",x"00300000",x"03DC00A0",x"037E000C",x"C57DFFFC",x"82003E98",x"07DC00A0",x"C05C0094",x"22640220",x"C09C0090",x"D4286000",x"8200D1FC",x"C4FC0090",x"C49C0094",x"C17DFFFC",x"004C0000",x"00300000",x"03DC00A0",x"037E000C",x"C57DFFFC",x"82003CC4",x"07DC00A0",x"C05C0094",x"22640220",x"C09C0090",x"D4286000",x"06240001",x"8620D3D4",x"22420220",x"C07C008C",x"D0464000",x"C09C0088",x"C0A80004",x"C0C80000",x"C0E40004",x"03000001",x"82F0D2A0",x"03000002",x"82F0D268",x"C4BC0098",x"C43C009C",x"C17DFFFC",x"002C0000",x"03DC00A8",x"037E000C",x"C57DFFFC",x"8200400C",x"07DC00A8",x"C05C009C",x"22640220",x"C09C0098",x"D4286000",x"8200D29C",x"C4BC0098",x"C43C009C",x"C17DFFFC",x"002C0000",x"03DC00A8",x"037E000C",x"C57DFFFC",x"82003E98",x"07DC00A8",x"C05C009C",x"22640220",x"C09C0098",x"D4286000",x"8200D2D4",x"C4BC0098",x"C43C009C",x"C17DFFFC",x"002C0000",x"03DC00A8",x"037E000C",x"C57DFFFC",x"82003CC4",x"07DC00A8",x"C05C009C",x"22640220",x"C09C0098",x"D4286000",x"06240001",x"8620D3D0",x"22420220",x"C07C008C",x"D0464000",x"C07C0088",x"C0860004",x"C0A60000",x"C0C40004",x"02E00001",x"82CED378",x"02E00002",x"82CED340",x"C49C00A0",x"C43C00A4",x"C17DFFFC",x"002A0000",x"03DC00B0",x"037E000C",x"C57DFFFC",x"8200400C",x"07DC00B0",x"C05C00A4",x"22640220",x"C09C00A0",x"D4286000",x"8200D374",x"C49C00A0",x"C43C00A4",x"C17DFFFC",x"002A0000",x"03DC00B0",x"037E000C",x"C57DFFFC",x"82003E98",x"07DC00B0",x"C05C00A4",x"22640220",x"C09C00A0",x"D4286000",x"8200D3AC",x"C49C00A0",x"C43C00A4",x"C17DFFFC",x"002A0000",x"03DC00B0",x"037E000C",x"C57DFFFC",x"82003CC4",x"07DC00B0",x"C05C00A4",x"22640220",x"C09C00A0",x"D4286000",x"06440001",x"C03C0088",x"C17DFFFC",x"03DC00B0",x"037E000C",x"C57DFFFC",x"820042A4",x"07DC00B0",x"8200D3D0",x"8200D3D4",x"8200D3D8",x"02400075",x"C03C006C",x"C17DFFFC",x"03DC00B0",x"037E000C",x"C57DFFFC",x"8200BD10",x"07DC00B0",x"C03C0068",x"06220001",x"8620D758",x"22420220",x"C07C0000",x"D0464000",x"C08401DC",x"C0BC0008",x"C0AA0000",x"06AA0001",x"C43C00A8",x"C45C00AC",x"86A0D6E8",x"02C000C8",x"22EA0220",x"D0ECE000",x"C1080004",x"C1280000",x"C14E0004",x"02600001",x"C49C00B0",x"C4DC00B4",x"8346D4D4",x"02600002",x"8346D498",x"C51C00B8",x"C4BC00BC",x"C17DFFFC",x"004E0000",x"00320000",x"03DC00C8",x"037E000C",x"C57DFFFC",x"8200400C",x"07DC00C8",x"C05C00BC",x"22640220",x"C09C00B8",x"D4286000",x"8200D4D0",x"C51C00B8",x"C4BC00BC",x"C17DFFFC",x"004E0000",x"00320000",x"03DC00C8",x"037E000C",x"C57DFFFC",x"82003E98",x"07DC00C8",x"C05C00BC",x"22640220",x"C09C00B8",x"D4286000",x"8200D50C",x"C51C00B8",x"C4BC00BC",x"C17DFFFC",x"004E0000",x"00320000",x"03DC00C8",x"037E000C",x"C57DFFFC",x"82003CC4",x"07DC00C8",x"C05C00BC",x"22640220",x"C09C00B8",x"D4286000",x"06240001",x"8620D6E4",x"22420220",x"C07C00B4",x"D0464000",x"C09C00B0",x"C0A80004",x"C0C80000",x"C0E40004",x"03000001",x"82F0D5B0",x"03000002",x"82F0D578",x"C4BC00C0",x"C43C00C4",x"C17DFFFC",x"002C0000",x"03DC00D0",x"037E000C",x"C57DFFFC",x"8200400C",x"07DC00D0",x"C05C00C4",x"22640220",x"C09C00C0",x"D4286000",x"8200D5AC",x"C4BC00C0",x"C43C00C4",x"C17DFFFC",x"002C0000",x"03DC00D0",x"037E000C",x"C57DFFFC",x"82003E98",x"07DC00D0",x"C05C00C4",x"22640220",x"C09C00C0",x"D4286000",x"8200D5E4",x"C4BC00C0",x"C43C00C4",x"C17DFFFC",x"002C0000",x"03DC00D0",x"037E000C",x"C57DFFFC",x"82003CC4",x"07DC00D0",x"C05C00C4",x"22640220",x"C09C00C0",x"D4286000",x"06240001",x"8620D6E0",x"22420220",x"C07C00B4",x"D0464000",x"C07C00B0",x"C0860004",x"C0A60000",x"C0C40004",x"02E00001",x"82CED688",x"02E00002",x"82CED650",x"C49C00C8",x"C43C00CC",x"C17DFFFC",x"002A0000",x"03DC00D8",x"037E000C",x"C57DFFFC",x"8200400C",x"07DC00D8",x"C05C00CC",x"22640220",x"C09C00C8",x"D4286000",x"8200D684",x"C49C00C8",x"C43C00CC",x"C17DFFFC",x"002A0000",x"03DC00D8",x"037E000C",x"C57DFFFC",x"82003E98",x"07DC00D8",x"C05C00CC",x"22640220",x"C09C00C8",x"D4286000",x"8200D6BC",x"C49C00C8",x"C43C00CC",x"C17DFFFC",x"002A0000",x"03DC00D8",x"037E000C",x"C57DFFFC",x"82003CC4",x"07DC00D8",x"C05C00CC",x"22640220",x"C09C00C8",x"D4286000",x"06440001",x"C03C00B0",x"C17DFFFC",x"03DC00D8",x"037E000C",x"C57DFFFC",x"820042A4",x"07DC00D8",x"8200D6E0",x"8200D6E4",x"8200D6E8",x"02400076",x"C03C00AC",x"C17DFFFC",x"03DC00D8",x"037E000C",x"C57DFFFC",x"8200BD10",x"07DC00D8",x"C03C00A8",x"06220001",x"8620D754",x"22420220",x"C07C0000",x"D0464000",x"02600077",x"C43C00D0",x"C17DFFFC",x"00240000",x"00460000",x"03DC00DC",x"037E000C",x"C57DFFFC",x"8200BD10",x"07DC00DC",x"C03C00D0",x"06220001",x"8200C714",x"C1FDFFFC",x"C1FDFFFC",x"C1FDFFFC",x"C1FDFFFC",x"22220220",x"02600640",x"C0860000",x"C82000A8",x"C044001C",x"C8440000",x"44224000",x"024001D0",x"C8440000",x"44404000",x"C8640004",x"44606000",x"C8840008",x"44808000",x"02A20001",x"C8A40000",x"02C00003",x"40C00000",x"C47C0000",x"CC5C0008",x"CCDC0010",x"C45C0018",x"C43C001C",x"C49C0020",x"C4BC0024",x"CC3C0028",x"CC9C0030",x"CC7C0038",x"CCBC0040",x"C17DFFFC",x"002C0000",x"4020C000",x"03DC0050",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0050",x"00420000",x"022000C4",x"C0620000",x"C43C0048",x"C45C004C",x"C17DFFFC",x"00260000",x"03DC0058",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0058",x"005A0000",x"03BA0008",x"C4240004",x"C07C004C",x"C4640000",x"C83C0040",x"CC260000",x"C83C0038",x"CC260004",x"C85C0030",x"CC460008",x"C09C0048",x"C0A80000",x"06AA0001",x"C45C0050",x"86A0DB00",x"02C000C8",x"22EA0220",x"D0ECE000",x"C10E0004",x"03200001",x"C4DC0054",x"8312D904",x"03200002",x"8312D8C8",x"C43C0058",x"C4BC005C",x"C17DFFFC",x"004E0000",x"00260000",x"03DC0068",x"037E000C",x"C57DFFFC",x"8200400C",x"07DC0068",x"C05C005C",x"22640220",x"C09C0058",x"D4286000",x"8200D900",x"C43C0058",x"C4BC005C",x"C17DFFFC",x"004E0000",x"00260000",x"03DC0068",x"037E000C",x"C57DFFFC",x"82003E98",x"07DC0068",x"C05C005C",x"22640220",x"C09C0058",x"D4286000",x"8200D93C",x"C43C0058",x"C4BC005C",x"C17DFFFC",x"004E0000",x"00260000",x"03DC0068",x"037E000C",x"C57DFFFC",x"82003CC4",x"07DC0068",x"C05C005C",x"22640220",x"C09C0058",x"D4286000",x"06240001",x"8620DAFC",x"22420220",x"C07C0054",x"D0464000",x"C0A40004",x"02C00001",x"82ACD9D4",x"02C00002",x"82ACD99C",x"C0BC004C",x"C43C0060",x"C17DFFFC",x"002A0000",x"03DC006C",x"037E000C",x"C57DFFFC",x"8200400C",x"07DC006C",x"C05C0060",x"22640220",x"C09C0058",x"D4286000",x"8200D9D0",x"C0BC004C",x"C43C0060",x"C17DFFFC",x"002A0000",x"03DC006C",x"037E000C",x"C57DFFFC",x"82003E98",x"07DC006C",x"C05C0060",x"22640220",x"C09C0058",x"D4286000",x"8200DA08",x"C0BC004C",x"C43C0060",x"C17DFFFC",x"002A0000",x"03DC006C",x"037E000C",x"C57DFFFC",x"82003CC4",x"07DC006C",x"C05C0060",x"22640220",x"C09C0058",x"D4286000",x"06240001",x"8620DAF8",x"22420220",x"C07C0054",x"D0464000",x"C0640004",x"02A00001",x"826ADAA0",x"02A00002",x"826ADA68",x"C07C004C",x"C43C0064",x"C17DFFFC",x"00260000",x"03DC0070",x"037E000C",x"C57DFFFC",x"8200400C",x"07DC0070",x"C05C0064",x"22640220",x"C09C0058",x"D4286000",x"8200DA9C",x"C07C004C",x"C43C0064",x"C17DFFFC",x"00260000",x"03DC0070",x"037E000C",x"C57DFFFC",x"82003E98",x"07DC0070",x"C05C0064",x"22640220",x"C09C0058",x"D4286000",x"8200DAD4",x"C07C004C",x"C43C0064",x"C17DFFFC",x"00260000",x"03DC0070",x"037E000C",x"C57DFFFC",x"82003CC4",x"07DC0070",x"C05C0064",x"22640220",x"C09C0058",x"D4286000",x"06440001",x"C03C0050",x"C17DFFFC",x"03DC0070",x"037E000C",x"C57DFFFC",x"820042A4",x"07DC0070",x"8200DAF8",x"8200DAFC",x"8200DB00",x"02200370",x"005A0000",x"03BA000C",x"C83C0028",x"CC240008",x"C07C0050",x"C4640004",x"C07C0024",x"C4640000",x"C07C0020",x"22860220",x"D4428000",x"02460001",x"C09C001C",x"02A80002",x"C0DC0018",x"C84C0004",x"02E00003",x"C87C0010",x"C43C0068",x"C45C006C",x"C4BC0070",x"CC5C0078",x"C17DFFFC",x"002E0000",x"40206000",x"03DC0088",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0088",x"00420000",x"C03C0048",x"C0620000",x"C45C0080",x"C17DFFFC",x"00260000",x"03DC008C",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC008C",x"005A0000",x"03BA0008",x"C4240004",x"C07C0080",x"C4640000",x"C83C0008",x"CC260000",x"C85C0078",x"CC460004",x"C85C0030",x"CC460008",x"C09C0048",x"C0A80000",x"06AA0001",x"C45C0084",x"86A0DE80",x"02C000C8",x"22EA0220",x"D0ECE000",x"C10E0004",x"03200001",x"C4DC0088",x"8312DC84",x"03200002",x"8312DC48",x"C43C008C",x"C4BC0090",x"C17DFFFC",x"004E0000",x"00260000",x"03DC009C",x"037E000C",x"C57DFFFC",x"8200400C",x"07DC009C",x"C05C0090",x"22640220",x"C09C008C",x"D4286000",x"8200DC80",x"C43C008C",x"C4BC0090",x"C17DFFFC",x"004E0000",x"00260000",x"03DC009C",x"037E000C",x"C57DFFFC",x"82003E98",x"07DC009C",x"C05C0090",x"22640220",x"C09C008C",x"D4286000",x"8200DCBC",x"C43C008C",x"C4BC0090",x"C17DFFFC",x"004E0000",x"00260000",x"03DC009C",x"037E000C",x"C57DFFFC",x"82003CC4",x"07DC009C",x"C05C0090",x"22640220",x"C09C008C",x"D4286000",x"06240001",x"8620DE7C",x"22420220",x"C07C0088",x"D0464000",x"C0A40004",x"02C00001",x"82ACDD54",x"02C00002",x"82ACDD1C",x"C0BC0080",x"C43C0094",x"C17DFFFC",x"002A0000",x"03DC00A0",x"037E000C",x"C57DFFFC",x"8200400C",x"07DC00A0",x"C05C0094",x"22640220",x"C09C008C",x"D4286000",x"8200DD50",x"C0BC0080",x"C43C0094",x"C17DFFFC",x"002A0000",x"03DC00A0",x"037E000C",x"C57DFFFC",x"82003E98",x"07DC00A0",x"C05C0094",x"22640220",x"C09C008C",x"D4286000",x"8200DD88",x"C0BC0080",x"C43C0094",x"C17DFFFC",x"002A0000",x"03DC00A0",x"037E000C",x"C57DFFFC",x"82003CC4",x"07DC00A0",x"C05C0094",x"22640220",x"C09C008C",x"D4286000",x"06240001",x"8620DE78",x"22420220",x"C07C0088",x"D0464000",x"C0640004",x"02A00001",x"826ADE20",x"02A00002",x"826ADDE8",x"C07C0080",x"C43C0098",x"C17DFFFC",x"00260000",x"03DC00A4",x"037E000C",x"C57DFFFC",x"8200400C",x"07DC00A4",x"C05C0098",x"22640220",x"C09C008C",x"D4286000",x"8200DE1C",x"C07C0080",x"C43C0098",x"C17DFFFC",x"00260000",x"03DC00A4",x"037E000C",x"C57DFFFC",x"82003E98",x"07DC00A4",x"C05C0098",x"22640220",x"C09C008C",x"D4286000",x"8200DE54",x"C07C0080",x"C43C0098",x"C17DFFFC",x"00260000",x"03DC00A4",x"037E000C",x"C57DFFFC",x"82003CC4",x"07DC00A4",x"C05C0098",x"22640220",x"C09C008C",x"D4286000",x"06440001",x"C03C0084",x"C17DFFFC",x"03DC00A4",x"037E000C",x"C57DFFFC",x"820042A4",x"07DC00A4",x"8200DE78",x"8200DE7C",x"8200DE80",x"003A0000",x"03BA000C",x"C83C0028",x"CC220008",x"C05C0084",x"C4420004",x"C05C0070",x"C4420000",x"C05C006C",x"22440220",x"C07C0068",x"D4264000",x"C03C0020",x"02420002",x"C09C001C",x"02880003",x"C0BC0018",x"C84A0008",x"02A00003",x"C87C0010",x"C45C009C",x"C49C00A0",x"CC5C00A8",x"C17DFFFC",x"002A0000",x"40206000",x"03DC00B8",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC00B8",x"00420000",x"C03C0048",x"C0620000",x"C45C00B0",x"C17DFFFC",x"00260000",x"03DC00BC",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC00BC",x"005A0000",x"03BA0008",x"C4240004",x"C07C00B0",x"C4640000",x"C83C0008",x"CC260000",x"C83C0038",x"CC260004",x"C83C00A8",x"CC260008",x"C09C0048",x"C0880000",x"06880001",x"C45C00B4",x"8680E200",x"02A000C8",x"22C80220",x"D0CAC000",x"C0EC0004",x"03000001",x"C4BC00B8",x"82F0E004",x"03000002",x"82F0DFC8",x"C43C00BC",x"C49C00C0",x"C17DFFFC",x"004C0000",x"00260000",x"03DC00CC",x"037E000C",x"C57DFFFC",x"8200400C",x"07DC00CC",x"C05C00C0",x"22640220",x"C09C00BC",x"D4286000",x"8200E000",x"C43C00BC",x"C49C00C0",x"C17DFFFC",x"004C0000",x"00260000",x"03DC00CC",x"037E000C",x"C57DFFFC",x"82003E98",x"07DC00CC",x"C05C00C0",x"22640220",x"C09C00BC",x"D4286000",x"8200E03C",x"C43C00BC",x"C49C00C0",x"C17DFFFC",x"004C0000",x"00260000",x"03DC00CC",x"037E000C",x"C57DFFFC",x"82003CC4",x"07DC00CC",x"C05C00C0",x"22640220",x"C09C00BC",x"D4286000",x"06240001",x"8620E1FC",x"22420220",x"C07C00B8",x"D0464000",x"C0A40004",x"02C00001",x"82ACE0D4",x"02C00002",x"82ACE09C",x"C0BC00B0",x"C43C00C4",x"C17DFFFC",x"002A0000",x"03DC00D0",x"037E000C",x"C57DFFFC",x"8200400C",x"07DC00D0",x"C05C00C4",x"22640220",x"C09C00BC",x"D4286000",x"8200E0D0",x"C0BC00B0",x"C43C00C4",x"C17DFFFC",x"002A0000",x"03DC00D0",x"037E000C",x"C57DFFFC",x"82003E98",x"07DC00D0",x"C05C00C4",x"22640220",x"C09C00BC",x"D4286000",x"8200E108",x"C0BC00B0",x"C43C00C4",x"C17DFFFC",x"002A0000",x"03DC00D0",x"037E000C",x"C57DFFFC",x"82003CC4",x"07DC00D0",x"C05C00C4",x"22640220",x"C09C00BC",x"D4286000",x"06240001",x"8620E1F8",x"22420220",x"C07C00B8",x"D0464000",x"C0640004",x"02A00001",x"826AE1A0",x"02A00002",x"826AE168",x"C07C00B0",x"C43C00C8",x"C17DFFFC",x"00260000",x"03DC00D4",x"037E000C",x"C57DFFFC",x"8200400C",x"07DC00D4",x"C05C00C8",x"22640220",x"C09C00BC",x"D4286000",x"8200E19C",x"C07C00B0",x"C43C00C8",x"C17DFFFC",x"00260000",x"03DC00D4",x"037E000C",x"C57DFFFC",x"82003E98",x"07DC00D4",x"C05C00C8",x"22640220",x"C09C00BC",x"D4286000",x"8200E1D4",x"C07C00B0",x"C43C00C8",x"C17DFFFC",x"00260000",x"03DC00D4",x"037E000C",x"C57DFFFC",x"82003CC4",x"07DC00D4",x"C05C00C8",x"22640220",x"C09C00BC",x"D4286000",x"06440001",x"C03C00B4",x"C17DFFFC",x"03DC00D4",x"037E000C",x"C57DFFFC",x"820042A4",x"07DC00D4",x"8200E1F8",x"8200E1FC",x"8200E200",x"003A0000",x"03BA000C",x"C83C0028",x"CC220008",x"C05C00B4",x"C4420004",x"C05C00A0",x"C4420000",x"C05C009C",x"22440220",x"C07C0068",x"D4264000",x"C03C0020",x"02220003",x"C05C0000",x"C4240000",x"C1FDFFFC",x"22220220",x"02220001",x"02600640",x"C0860000",x"C82000A8",x"C0A4001C",x"C84A0000",x"44224000",x"02A001D0",x"C0C40010",x"C84A0000",x"C86C0000",x"48446000",x"C86A0004",x"C88C0004",x"48668000",x"40446000",x"C86A0008",x"C88C0008",x"48668000",x"40446000",x"C8600080",x"C0C40010",x"C88C0000",x"48868000",x"48884000",x"C8AA0000",x"4488A000",x"C0C40010",x"C8AC0004",x"48A6A000",x"48AA4000",x"C8CA0004",x"44AAC000",x"C0440010",x"C8C40008",x"4866C000",x"48464000",x"C86A0008",x"44446000",x"02400003",x"40600000",x"C47C0000",x"C49C0004",x"C43C0008",x"CC3C0010",x"CC5C0018",x"CCBC0020",x"CC9C0028",x"C17DFFFC",x"00240000",x"40206000",x"03DC0038",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0038",x"00420000",x"022000C4",x"C0620000",x"C43C0030",x"C45C0034",x"C17DFFFC",x"00260000",x"03DC0040",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0040",x"005A0000",x"03BA0008",x"C4240004",x"C07C0034",x"C4640000",x"C83C0028",x"CC260000",x"C83C0020",x"CC260004",x"C83C0018",x"CC260008",x"C09C0030",x"C0880000",x"06880001",x"C45C0038",x"8680E630",x"02A000C8",x"22C80220",x"D0CAC000",x"C0EC0004",x"03000001",x"C4BC003C",x"82F0E434",x"03000002",x"82F0E3F8",x"C43C0040",x"C49C0044",x"C17DFFFC",x"004C0000",x"00260000",x"03DC0050",x"037E000C",x"C57DFFFC",x"8200400C",x"07DC0050",x"C05C0044",x"22640220",x"C09C0040",x"D4286000",x"8200E430",x"C43C0040",x"C49C0044",x"C17DFFFC",x"004C0000",x"00260000",x"03DC0050",x"037E000C",x"C57DFFFC",x"82003E98",x"07DC0050",x"C05C0044",x"22640220",x"C09C0040",x"D4286000",x"8200E46C",x"C43C0040",x"C49C0044",x"C17DFFFC",x"004C0000",x"00260000",x"03DC0050",x"037E000C",x"C57DFFFC",x"82003CC4",x"07DC0050",x"C05C0044",x"22640220",x"C09C0040",x"D4286000",x"06240001",x"8620E62C",x"22420220",x"C07C003C",x"D0464000",x"C0A40004",x"02C00001",x"82ACE504",x"02C00002",x"82ACE4CC",x"C0BC0034",x"C43C0048",x"C17DFFFC",x"002A0000",x"03DC0054",x"037E000C",x"C57DFFFC",x"8200400C",x"07DC0054",x"C05C0048",x"22640220",x"C09C0040",x"D4286000",x"8200E500",x"C0BC0034",x"C43C0048",x"C17DFFFC",x"002A0000",x"03DC0054",x"037E000C",x"C57DFFFC",x"82003E98",x"07DC0054",x"C05C0048",x"22640220",x"C09C0040",x"D4286000",x"8200E538",x"C0BC0034",x"C43C0048",x"C17DFFFC",x"002A0000",x"03DC0054",x"037E000C",x"C57DFFFC",x"82003CC4",x"07DC0054",x"C05C0048",x"22640220",x"C09C0040",x"D4286000",x"06240001",x"8620E628",x"22420220",x"C07C003C",x"D0464000",x"C0640004",x"02A00001",x"826AE5D0",x"02A00002",x"826AE598",x"C07C0034",x"C43C004C",x"C17DFFFC",x"00260000",x"03DC0058",x"037E000C",x"C57DFFFC",x"8200400C",x"07DC0058",x"C05C004C",x"22640220",x"C09C0040",x"D4286000",x"8200E5CC",x"C07C0034",x"C43C004C",x"C17DFFFC",x"00260000",x"03DC0058",x"037E000C",x"C57DFFFC",x"82003E98",x"07DC0058",x"C05C004C",x"22640220",x"C09C0040",x"D4286000",x"8200E604",x"C07C0034",x"C43C004C",x"C17DFFFC",x"00260000",x"03DC0058",x"037E000C",x"C57DFFFC",x"82003CC4",x"07DC0058",x"C05C004C",x"22640220",x"C09C0040",x"D4286000",x"06440001",x"C03C0038",x"C17DFFFC",x"03DC0058",x"037E000C",x"C57DFFFC",x"820042A4",x"07DC0058",x"8200E628",x"8200E62C",x"8200E630",x"02200370",x"005A0000",x"03BA000C",x"C83C0010",x"CC240008",x"C07C0038",x"C4640004",x"C07C0008",x"C4640000",x"C07C0004",x"22860220",x"D4428000",x"02260001",x"C05C0000",x"C4240000",x"C1FDFFFC",x"026002F8",x"C4260000",x"C4460004",x"02800300",x"22A201A0",x"C4A80000",x"224401A0",x"C4480004",x"02400308",x"C8200004",x"58420000",x"C47C0000",x"C45C0004",x"CC3C0008",x"C17DFFFC",x"40204000",x"03DC0018",x"037E000C",x"C57DFFFC",x"82000844",x"07DC0018",x"C85C0008",x"48242000",x"C03C0004",x"CC220000",x"C03C0000",x"C0420000",x"C45C0010",x"C17DFFFC",x"03DC001C",x"037E000C",x"C57DFFFC",x"8200A47C",x"07DC001C",x"00420000",x"C03C0010",x"C17DFFFC",x"03DC001C",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC001C",x"C05C0000",x"C0640000",x"06660002",x"C17DFFFC",x"00460000",x"03DC001C",x"037E000C",x"C57DFFFC",x"8200A914",x"07DC001C",x"C05C0000",x"C0640000",x"C43C0014",x"C47C0018",x"C17DFFFC",x"03DC0024",x"037E000C",x"C57DFFFC",x"8200A47C",x"07DC0024",x"00420000",x"C03C0018",x"C17DFFFC",x"03DC0024",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0024",x"C05C0000",x"C0640000",x"06660002",x"C17DFFFC",x"00460000",x"03DC0024",x"037E000C",x"C57DFFFC",x"8200A914",x"07DC0024",x"C05C0000",x"C0640000",x"C43C001C",x"C47C0020",x"C17DFFFC",x"03DC002C",x"037E000C",x"C57DFFFC",x"8200A47C",x"07DC002C",x"00420000",x"C03C0020",x"C17DFFFC",x"03DC002C",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC002C",x"C05C0000",x"C0640000",x"06660002",x"C17DFFFC",x"00460000",x"03DC002C",x"037E000C",x"C57DFFFC",x"8200A914",x"07DC002C",x"C43C0024",x"C17DFFFC",x"03DC0030",x"037E000C",x"C57DFFFC",x"820016D4",x"07DC0030",x"C17DFFFC",x"03DC0030",x"037E000C",x"C57DFFFC",x"82001AB8",x"07DC0030",x"02200000",x"C43C0028",x"C17DFFFC",x"03DC0034",x"037E000C",x"C57DFFFC",x"82002384",x"07DC0034",x"8220E898",x"02200001",x"C17DFFFC",x"03DC0034",x"037E000C",x"C57DFFFC",x"82002930",x"07DC0034",x"8200E8A4",x"022000C4",x"C05C0028",x"C4420000",x"C17DFFFC",x"03DC0034",x"037E000C",x"C57DFFFC",x"82000794",x"07DC0034",x"0240FFFF",x"8224E8F4",x"02400001",x"C43C002C",x"C17DFFFC",x"00240000",x"03DC0038",x"037E000C",x"C57DFFFC",x"82002A44",x"07DC0038",x"C05C002C",x"C4420000",x"8200E914",x"02200001",x"0240FFFF",x"C17DFFFC",x"03DC0038",x"037E000C",x"C57DFFFC",x"8200081C",x"07DC0038",x"C0420000",x"0260FFFF",x"8246E980",x"024001E0",x"C4240000",x"02200000",x"C45C0030",x"C17DFFFC",x"03DC003C",x"037E000C",x"C57DFFFC",x"82002A44",x"07DC003C",x"C0420000",x"0260FFFF",x"8246E97C",x"C05C0030",x"C4240004",x"02200002",x"C17DFFFC",x"03DC003C",x"037E000C",x"C57DFFFC",x"82002E74",x"07DC003C",x"8200E97C",x"8200E980",x"022002A8",x"02400000",x"C43C0034",x"C17DFFFC",x"00240000",x"03DC0040",x"037E000C",x"C57DFFFC",x"82002BEC",x"07DC0040",x"C05C0034",x"C4240000",x"02200050",x"C17DFFFC",x"03DC0040",x"037E000C",x"C57DFFFC",x"8200078C",x"07DC0040",x"02200036",x"C17DFFFC",x"03DC0040",x"037E000C",x"C57DFFFC",x"8200078C",x"07DC0040",x"0220000A",x"C17DFFFC",x"03DC0040",x"037E000C",x"C57DFFFC",x"8200078C",x"07DC0040",x"02200031",x"C17DFFFC",x"03DC0040",x"037E000C",x"C57DFFFC",x"8200078C",x"07DC0040",x"02200032",x"C17DFFFC",x"03DC0040",x"037E000C",x"C57DFFFC",x"8200078C",x"07DC0040",x"02200038",x"C17DFFFC",x"03DC0040",x"037E000C",x"C57DFFFC",x"8200078C",x"07DC0040",x"02200020",x"C17DFFFC",x"03DC0040",x"037E000C",x"C57DFFFC",x"8200078C",x"07DC0040",x"02200031",x"C17DFFFC",x"03DC0040",x"037E000C",x"C57DFFFC",x"8200078C",x"07DC0040",x"02200032",x"C17DFFFC",x"03DC0040",x"037E000C",x"C57DFFFC",x"8200078C",x"07DC0040",x"02200038",x"C17DFFFC",x"03DC0040",x"037E000C",x"C57DFFFC",x"8200078C",x"07DC0040",x"0220000A",x"C17DFFFC",x"03DC0040",x"037E000C",x"C57DFFFC",x"8200078C",x"07DC0040",x"02200032",x"C17DFFFC",x"03DC0040",x"037E000C",x"C57DFFFC",x"8200078C",x"07DC0040",x"02200035",x"C17DFFFC",x"03DC0040",x"037E000C",x"C57DFFFC",x"8200078C",x"07DC0040",x"02200035",x"C17DFFFC",x"03DC0040",x"037E000C",x"C57DFFFC",x"8200078C",x"07DC0040",x"0220000A",x"C17DFFFC",x"03DC0040",x"037E000C",x"C57DFFFC",x"8200078C",x"07DC0040",x"02200004",x"C17DFFFC",x"03DC0040",x"037E000C",x"C57DFFFC",x"8200B92C",x"07DC0040",x"02200009",x"02400000",x"02600000",x"C17DFFFC",x"03DC0040",x"037E000C",x"C57DFFFC",x"8200B574",x"07DC0040",x"02200354",x"C0420010",x"C06401DC",x"028000C4",x"C0A80000",x"06AA0001",x"C49C0038",x"C43C003C",x"C45C0040",x"86A0EE78",x"02C000C8",x"22EA0220",x"D0ECE000",x"C1060004",x"C1260000",x"C14E0004",x"02800001",x"C47C0044",x"C4DC0048",x"8348EC64",x"02800002",x"8348EC28",x"C51C004C",x"C4BC0050",x"C17DFFFC",x"004E0000",x"00320000",x"03DC005C",x"037E000C",x"C57DFFFC",x"8200400C",x"07DC005C",x"C05C0050",x"22640220",x"C09C004C",x"D4286000",x"8200EC60",x"C51C004C",x"C4BC0050",x"C17DFFFC",x"004E0000",x"00320000",x"03DC005C",x"037E000C",x"C57DFFFC",x"82003E98",x"07DC005C",x"C05C0050",x"22640220",x"C09C004C",x"D4286000",x"8200EC9C",x"C51C004C",x"C4BC0050",x"C17DFFFC",x"004E0000",x"00320000",x"03DC005C",x"037E000C",x"C57DFFFC",x"82003CC4",x"07DC005C",x"C05C0050",x"22640220",x"C09C004C",x"D4286000",x"06240001",x"8620EE74",x"22420220",x"C07C0048",x"D0464000",x"C09C0044",x"C0A80004",x"C0C80000",x"C0E40004",x"03000001",x"82F0ED40",x"03000002",x"82F0ED08",x"C4BC0054",x"C43C0058",x"C17DFFFC",x"002C0000",x"03DC0064",x"037E000C",x"C57DFFFC",x"8200400C",x"07DC0064",x"C05C0058",x"22640220",x"C09C0054",x"D4286000",x"8200ED3C",x"C4BC0054",x"C43C0058",x"C17DFFFC",x"002C0000",x"03DC0064",x"037E000C",x"C57DFFFC",x"82003E98",x"07DC0064",x"C05C0058",x"22640220",x"C09C0054",x"D4286000",x"8200ED74",x"C4BC0054",x"C43C0058",x"C17DFFFC",x"002C0000",x"03DC0064",x"037E000C",x"C57DFFFC",x"82003CC4",x"07DC0064",x"C05C0058",x"22640220",x"C09C0054",x"D4286000",x"06240001",x"8620EE70",x"22420220",x"C07C0048",x"D0464000",x"C07C0044",x"C0860004",x"C0A60000",x"C0C40004",x"02E00001",x"82CEEE18",x"02E00002",x"82CEEDE0",x"C49C005C",x"C43C0060",x"C17DFFFC",x"002A0000",x"03DC006C",x"037E000C",x"C57DFFFC",x"8200400C",x"07DC006C",x"C05C0060",x"22640220",x"C09C005C",x"D4286000",x"8200EE14",x"C49C005C",x"C43C0060",x"C17DFFFC",x"002A0000",x"03DC006C",x"037E000C",x"C57DFFFC",x"82003E98",x"07DC006C",x"C05C0060",x"22640220",x"C09C005C",x"D4286000",x"8200EE4C",x"C49C005C",x"C43C0060",x"C17DFFFC",x"002A0000",x"03DC006C",x"037E000C",x"C57DFFFC",x"82003CC4",x"07DC006C",x"C05C0060",x"22640220",x"C09C005C",x"D4286000",x"06440001",x"C03C0044",x"C17DFFFC",x"03DC006C",x"037E000C",x"C57DFFFC",x"820042A4",x"07DC006C",x"8200EE70",x"8200EE74",x"8200EE78",x"02400076",x"C03C0040",x"C17DFFFC",x"03DC006C",x"037E000C",x"C57DFFFC",x"8200BD10",x"07DC006C",x"C03C003C",x"C022000C",x"02400077",x"C17DFFFC",x"03DC006C",x"037E000C",x"C57DFFFC",x"8200BD10",x"07DC006C",x"02200002",x"C17DFFFC",x"03DC006C",x"037E000C",x"C57DFFFC",x"8200C714",x"07DC006C",x"02200368",x"C0420000",x"026001D0",x"C8260000",x"CC240000",x"C8260004",x"CC240004",x"C8260008",x"CC240008",x"C05C0038",x"C0640000",x"06660001",x"8660F0EC",x"028000C8",x"22A60220",x"D0A8A000",x"C0C20004",x"C0E20000",x"C10A0004",x"03200001",x"C43C0064",x"C49C0068",x"8312EFB4",x"03200002",x"8312EF78",x"C4DC006C",x"C47C0070",x"C17DFFFC",x"004A0000",x"002E0000",x"03DC007C",x"037E000C",x"C57DFFFC",x"8200400C",x"07DC007C",x"C05C0070",x"22640220",x"C09C006C",x"D4286000",x"8200EFB0",x"C4DC006C",x"C47C0070",x"C17DFFFC",x"004A0000",x"002E0000",x"03DC007C",x"037E000C",x"C57DFFFC",x"82003E98",x"07DC007C",x"C05C0070",x"22640220",x"C09C006C",x"D4286000",x"8200EFEC",x"C4DC006C",x"C47C0070",x"C17DFFFC",x"004A0000",x"002E0000",x"03DC007C",x"037E000C",x"C57DFFFC",x"82003CC4",x"07DC007C",x"C05C0070",x"22640220",x"C09C006C",x"D4286000",x"06240001",x"8620F0E8",x"22420220",x"C07C0068",x"D0464000",x"C07C0064",x"C0860004",x"C0A60000",x"C0C40004",x"02E00001",x"82CEF090",x"02E00002",x"82CEF058",x"C49C0074",x"C43C0078",x"C17DFFFC",x"002A0000",x"03DC0084",x"037E000C",x"C57DFFFC",x"8200400C",x"07DC0084",x"C05C0078",x"22640220",x"C09C0074",x"D4286000",x"8200F08C",x"C49C0074",x"C43C0078",x"C17DFFFC",x"002A0000",x"03DC0084",x"037E000C",x"C57DFFFC",x"82003E98",x"07DC0084",x"C05C0078",x"22640220",x"C09C0074",x"D4286000",x"8200F0C4",x"C49C0074",x"C43C0078",x"C17DFFFC",x"002A0000",x"03DC0084",x"037E000C",x"C57DFFFC",x"82003CC4",x"07DC0084",x"C05C0078",x"22640220",x"C09C0074",x"D4286000",x"06440001",x"C03C0064",x"C17DFFFC",x"03DC0084",x"037E000C",x"C57DFFFC",x"820042A4",x"07DC0084",x"8200F0E8",x"8200F0EC",x"C03C0038",x"C0220000",x"06220001",x"8620F17C",x"024000C8",x"22620220",x"D0446000",x"C0640008",x"02800002",x"8268F118",x"8200F178",x"C064001C",x"C8260000",x"C84000A8",x"8E24F12C",x"8200F178",x"C0640004",x"02800001",x"8268F160",x"02800002",x"8268F144",x"8200F15C",x"C17DFFFC",x"03DC0084",x"037E000C",x"C57DFFFC",x"8200E244",x"07DC0084",x"8200F178",x"C17DFFFC",x"03DC0084",x"037E000C",x"C57DFFFC",x"8200D764",x"07DC0084",x"8200F17C",x"02400000",x"02600000",x"C03C001C",x"C17DFFFC",x"03DC0084",x"037E000C",x"C57DFFFC",x"82009C08",x"07DC0084",x"02400000",x"02600002",x"C03C0000",x"C0820004",x"8608F1B8",x"C1FDFFFC",x"C0220004",x"06220001",x"C45C007C",x"8602F1CC",x"8200F1F4",x"02200001",x"C09C0024",x"C17DFFFC",x"00420000",x"00280000",x"03DC0088",x"037E000C",x"C57DFFFC",x"82009C08",x"07DC0088",x"02200000",x"C05C007C",x"C07C0014",x"C09C001C",x"C0BC0024",x"C17DFFFC",x"03DC0088",x"037E000C",x"C57DFFFC",x"82009C7C",x"07DC0088",x"02200001",x"02A00004",x"C05C001C",x"C07C0024",x"C09C0014",x"C17DFFFC",x"03DC0088",x"037E000C",x"C57DFFFC",x"8200A164",x"07DC0088",x"C1FDFFFC",x"03DC0004",x"037E000C",x"C57DFFFC",x"82000644",x"07DC0004",x"02200080",x"02400080",x"C17DFFFC",x"03DC0008",x"037E000C",x"C57DFFFC",x"8200E670",x"07DC0008",x"02200000",x"8001E000",others => x"00000000");
  type cache_addr_array is array(16383 downto 0) of std_logic_vector(19 downto 0);
  signal cache_inst_addr : cache_addr_array := (others => x"FFFFF");
  signal cache_found : std_logic := '0';
begin
  with_alu: alu Port map (
      clk => clk,
      opc_alu => opccode_alu,
      reg_in_a => reg_in_a,
      reg_in_b => reg_in_b,
      reg_out => reg_out,
      shift_dir => shift_dir,
      shift_type => shift_type,
      shift_go => shift_go
    );
  with_compr: compr Port map (
      clk => clk,
      opc_compr => opccode_compr,
      reg_in_a => reg_in_a_compr,
      reg_in_b => reg_in_b_compr,
      cond_out => cond_out_compr
    );
  with_fpu: fpu_man Port map (
      clk => clk,
      opc_fpu => opccode_fpu,
      reg_in_a => reg_in_a_fpu,
      reg_in_b => reg_in_b_fpu,
      reg_out => reg_out_fpu
    );
  core_pro: process(clk)
    variable ftdcode : std_logic_vector(31 downto 0);
  begin
    if (rising_edge(clk)) and (execute_ok = '1') then
      -- state action one
      if state = x"00" then
        -- initialize groups
        if phase = "000" then
          --Phase Fetch
          --if waitwrite_from_parent = 0 then
            --if (rg(15)(31 downto 2)) < 110 then
            cache_found <= '1';
            --if cache_inst_addr(conv_integer(rg(15)(15 downto 2))) = (rg(15) (31 downto 12)) then
              -- cache match
            --  cache_found <= '1';
            --else
              -- cache mismatch
            --  cache_found <= '0';
            --  waitwriting <= '0';
            --  sram_go <= '1';
            --  sram_addr <= rg (15) (21 downto 2);
            --  sram_inst_type <= '0';
            --end if;
          --else
          --  waitwriting <= '1';
          --end if;
        end if;
        if phase = "010" then
          --Phase Decode and Load (Decode Side)
          --if waitwrite_from_parent = 0 then
            if cache_found = '1' then
              ftdcode := cache_inst(conv_integer(rg(15)(15 downto 2)));
            else
              ftdcode := sram_read;
              -- update cache
              cache_inst(conv_integer(rg(15)(15 downto 2))) <= sram_read;
              cache_inst_addr(conv_integer(rg(15)(15 downto 2))) <= (rg(15) (31 downto 12));
            end if;
            --ftdcode := sram_read;
          --else
            --nop
          --  ftdcode := x"FFFFFFFF";
          --end if;
          if (waitwrite_from_parent > 0) and (ftdcode(31 downto 25) = "1110001") then
            --write wait
            ftdcode := x"FFFFFFFF";
          end if;
          --Phase Decode and Load (Load Side)
          -- ALU
          if ftdcode(31 downto 30) = "00" then
            --set source A
            loaded_srca <= rg (conv_integer (ftdcode(20 downto 17)));
            --set source B
            if (ftdcode(31 downto 25) = "0000001") or (ftdcode(31 downto 25) = "0000011") or (ftdcode(31 downto 25) = "0010001") then
              --immediate
              if ftdcode(31 downto 25) = "0010001" then
                loaded_srcb <= x"000000" & "000" & ftdcode(12 downto 8);
              else
                if ftdcode(16) = '1' then
                  -- high
                  loaded_srcb <= ftdcode(15 downto 0)&"0000000000000000";
                else
                  -- low
                  if ftdcode(15) = '1' then
                    loaded_srcb <= "1111111111111111"&ftdcode(15 downto 0);
                  else
                    loaded_srcb <= "0000000000000000"&ftdcode(15 downto 0);
                  end if;
                end if;
              end if;
            else
              loaded_srcb <= rg (conv_integer (ftdcode(16 downto 13)));
            end if;
          end if;
          --FPU
          if ftdcode(31 downto 30) = "01" then
            --set source A
            if ftdcode(31 downto 25) = "0101100" then
              -- itof
              loaded_srca <= rg (conv_integer (ftdcode(20 downto 17)));
            else
              -- otherwise
              loaded_srca <= fp (conv_integer(ftdcode(20 downto 17)));
            end if;
            --set source B
            loaded_srcb <= fp (conv_integer (ftdcode(16 downto 13)));
          end if;
          --Branch
          if ftdcode(31 downto 30) = "10" then
            if ftdcode(31 downto 27) = "10001" then
              --float
              --set source A
              loaded_srca <= fp (conv_integer (ftdcode(24 downto 21)));
              --set source B
              loaded_srcb <= fp (conv_integer (ftdcode(20 downto 17)));
            else
              --integer
              --set source A
              loaded_srca <= rg (conv_integer(ftdcode(24 downto 21)));
              --set source B
              loaded_srcb <= rg (conv_integer (ftdcode(20 downto 17)));
            end if;
            --set newpc
            loaded_newpc <= rg (conv_integer(ftdcode(16 downto 13)));
          end if;
        end if;
        if phase = "011" then
          --Phase EXEC
          --ALU
          if ftdcode(31 downto 30) = "00" then
            opccode_alu <= ftdcode(31 downto 25);
            reg_in_a <= loaded_srca;
            reg_in_b <= loaded_srcb;
            if ftdcode(31 downto 29) = "001" then
              shift_dir <= ftdcode(7);
              shift_type <= ftdcode(6 downto 5);
              shift_go <= '1';
            end if;
          end if;
          --FPU
          if ftdcode(31 downto 30) = "01" then
            opccode_fpu <= ftdcode(31 downto 25);
            reg_in_a_fpu <= loaded_srca;
            reg_in_b_fpu <= loaded_srcb;
          end if;
          --Branch
          if ftdcode(31 downto 30) = "10" then
            if ftdcode(31 downto 27) = "10001" then
              opccode_fpu <= ftdcode(31 downto 25);
              reg_in_a_fpu <= loaded_srca;
              reg_in_b_fpu <= loaded_srcb;
            else
              opccode_compr <= ftdcode(31 downto 25);
              reg_in_a_compr <= loaded_srca;
              reg_in_b_compr <= loaded_srcb;
            end if;
            --Calculate next PC if branch condition is true
            opccode_alu <= "0000000";
            if ftdcode(25 downto 25) = "1" then
              -- branch imm type
              reg_in_a <= rg (0);
              reg_in_b <= x"000" & "000" & ftdcode(16 downto 0);
            else
              -- branch reg+imm type
              reg_in_a <= loaded_newpc;
              if ftdcode(12) = '1' then
                reg_in_b <= x"FFFF" & "111" & ftdcode(12 downto 0);
              else
                reg_in_b <= x"0000" & "000" & ftdcode(12 downto 0);
              end if;
            end if;
          end if;
          --MEMORY
          if (ftdcode(31 downto 25) = "1100000") or (ftdcode(31 downto 25) = "1101000") or (ftdcode(31 downto 25) = "1100100") or (ftdcode(31 downto 25) = "1101100") then
            --load, loadr, fload, floadr
            --calculate address
            --register A
            reg_in_a <= rg (conv_integer (ftdcode(20 downto 17)));
            --register B
            if ftdcode(28) = '0' then
              --load, fload
              if ftdcode(16) = '1' then
                reg_in_b <= x"FFF" & "111" & ftdcode(16 downto 0);
              else
                reg_in_b <= x"000" & "000" & ftdcode(16 downto 0);
              end if;
            else
              --loadr, floadr
              reg_in_b <= rg (conv_integer(ftdcode(16 downto 13)));
            end if;
            opccode_alu <= "0000000";
          end if;
          if (ftdcode(31 downto 25) = "1100010") or (ftdcode(31 downto 25) = "1101010") or (ftdcode(31 downto 25) = "1100110") or (ftdcode(31 downto 25) = "1101110") then
            --store, storer, fstore, fstorer
            reg_in_a <= rg (conv_integer(ftdcode(20 downto 17)));
            --register B
            if ftdcode(28) = '0' then
              --store, fstore
              if ftdcode(16) = '1' then
                reg_in_b <= x"FFF" & "111" & ftdcode(16 downto 0);
              else
                reg_in_b <= x"000" & "000" & ftdcode(16 downto 0);
              end if;
            else
              --storer, fstorer
              reg_in_b <= rg (conv_integer(ftdcode(16 downto 13)));
            end if;
            opccode_alu <= "0000000";
          end if;
          if ftdcode(31 downto 25) = "1110001" then
            -- write
            if ftdcode(24 downto 21) /= x"0" then
              debug_otpt <= rg (conv_integer(ftdcode(24 downto 21))) (7 downto 0);
            end if;
            debug_otpt_signal <= '1';
          else
            --if ftdcode(31 downto 20) = x"FFD" then
            ---- Debug Output
            --  if ftdcode(3 downto 0) = x"1" then
            --    debug_otpt <= rg(1) (7 downto 0);
            --  end if;
            --  if ftdcode(3 downto 0) = x"2" then
            --    debug_otpt <= rg(2) (7 downto 0);
            --  end if;
            --  if ftdcode(3 downto 0) = x"3" then
            --    debug_otpt <= rg(3) (7 downto 0);
            --  end if;
            --  debug_otpt_signal <= '1';
            --else
              debug_otpt_signal <= '0';
            --end if;
          end if;
          -- Debug NOP(all FFFFFFF case doesn't update PC)
        else
          -- the case state = 0 ^ phase != 100
          debug_otpt_signal <= '0';
        end if;
        if phase = "100" then
          --MEMORY
          --Phase Store
          --ALU
          if ftdcode(31 downto 30) = "00" then
            if ftdcode(24 downto 21) /= x"0" then
              rg (conv_integer(ftdcode(24 downto 21))) <= reg_out;
            end if;
          end if;
          --FPU
          if ftdcode(31 downto 30) = "01" then
            if ftdcode(31 downto 25) = "0101010" then
              --ftoi
              if ftdcode(24 downto 21) /= x"0" then
                rg (conv_integer(ftdcode(24 downto 21))) <= reg_out_fpu;
              end if;
            else
              if ftdcode(24 downto 21) /= x"0" then
                fp (conv_integer (ftdcode(24 downto 21))) <= reg_out_fpu;
              end if;
            end if;
          end if;
          if (ftdcode(31 downto 25) = "1100000") or (ftdcode(31 downto 25) = "1101000") then
            --load,loadr(integer)
            if ftdcode(24 downto 21) /= x"0" then
              if reg_out(21 downto 2) < 15522 then
                rg (conv_integer (ftdcode(24 downto 21))) <= cache_inst (conv_integer (reg_out(21 downto 2)));
              else
                rg (conv_integer (ftdcode(24 downto 21))) <= sram_read;
              end if;
            end if;
          end if;
          if (ftdcode(31 downto 25) = "1100100") or (ftdcode(31 downto 25) = "1101100") then
            --fload,floadr(float)
            if ftdcode(24 downto 21) /= x"0" then
              if reg_out(21 downto 2) < 15522 then
                fp (conv_integer (ftdcode(24 downto 21))) <= cache_inst (conv_integer (reg_out(21 downto 2)));
              else
                fp (conv_integer (ftdcode(24 downto 21))) <= sram_read;
              end if;
            end if;
          end if;
          if ftdcode(31 downto 25) = "1110000" then
            --read
            if ftdcode(24 downto 21) /= x"0" then
              rg (conv_integer(ftdcode(24 downto 21))) <= sram_read;
            end if;
            -- hp <= hp + 4
--            rg (13) <= rg (13) + 4;
          end if;
          --Update PC (Branch case)
          if ftdcode(31 downto 30) = "10" then
            --pc <= cond_new_pc;
            rg (15) <= cond_new_pc;
          else
            if ftdcode(31 downto 0) = x"FFFFFFFF" then
              -- added nop
            else
              -- The Case when update pc by ALU,load,loadr
              if ((ftdcode(31 downto 30) = "00") or (ftdcode(31 downto 25) = "0101010")) and (ftdcode(24 downto 21) = x"F") then
              else
                if ((ftdcode(31 downto 25) = "1100000") or (ftdcode(31 downto 25) = "1101000")) and (ftdcode(24 downto 21) = x"F") then
                else
                  --pc <= pc + 4;   
                  rg (15) <= rg (15) + 4;
                end if;
              end if;
            end if;
          end if;
        end if;
      else
        -- the case state != 0
        debug_otpt_signal <= '0';
      end if;
      if state = x"01" then
        sram_go <= '0';
        shift_go <= '0';
      end if;
      -- state action two
      if state = x"80" then
        if phase = "011" then
          --Phase EXEC
          if (ftdcode(31 downto 25) = "1100000") or (ftdcode(31 downto 25) = "1101000") or (ftdcode(31 downto 25) = "1100100") or (ftdcode(31 downto 25) = "1101100") then
            --load,loadr,fload,floadr
            sram_go <= '1';
            sram_addr <= reg_out(21 downto 2);
            sram_inst_type <= '0';
          end if;
          if (ftdcode(31 downto 25) = "1100010") or (ftdcode(31 downto 25) = "1101010") then
            --store,storer(integer)
            sram_go <= '1';
            sram_inst_type <= '1';
            sram_addr <= reg_out(21 downto 2);
            sram_write <= rg (conv_integer (ftdcode(24 downto 21)));
          end if;
          if (ftdcode(31 downto 25) = "1100110") or (ftdcode(31 downto 25) = "1101110") then
            --fstore,fstorer(float)
            sram_go <= '1';
            sram_inst_type <= '1';
            sram_addr <= reg_out(21 downto 2);
            sram_write <= fp (conv_integer (ftdcode(24 downto 21)));
          end if;
          if ftdcode(31 downto 25) = "1110000" then
            --read
--            sram_go <= '1';
              read_signal <= '1';
            -- sram_addr <= hp(21 downto 2);
--            sram_addr <= rg (13) (21 downto 2);
--            sram_inst_type <= '0';
          end if;
          -- pickup groups
          -- Update cond_new_pc
          if ftdcode(31 downto 27) = "10001" then
            if reg_out_fpu(0) = '1' then
              cond_new_pc <= reg_out;
            else
              -- cond_new_pc <= pc + 4;
              cond_new_pc <= rg (15) + 4;
            end if;            
          else
            if cond_out_compr = '1' then
              cond_new_pc <= reg_out;
            else
              -- cond_new_pc <= pc + 4;
              cond_new_pc <= rg (15) + 4;
            end if;
          end if;
        else
          sram_go <= '0';
        end if;
      end if;
      if state = x"81" then
        --reflesh
        sram_go <= '0';
        read_signal <= '0';
      end if;
      --if state = x"BB" then
      --  debug_otpt <= reg_out;
      --end if;
      if state = x"FF" then
        -- move to next phase
        phase <= phase + 1;
      end if;
      --state update
      if phase = "000" then
        -- Fetch
        if state = x"EA" then
          --skip
          state <= x"FF";
--          phase <= "010";
--          state <= x"00";
        elsif state = x"01" then
          --skip
          if (cache_found = '1') or (waitwriting = '1') then
            state <= x"FF";
--            phase <= "010";
--            state <= x"00";
          else
            state <= x"E0";
          end if;
        elsif state = x"FF" then
          phase <= "010";
          state <= x"00";
        else
          state <= state + 1;
        end if;
      end if;
      if phase = "010" then
        -- Load
        if state = x"01" then
          --skip
--          state <= x"FF";
          state <= x"00";
          phase <= phase + 1;
        else
          state <= state + 1;
        end if;
      end if;
      if phase = "011" then
        -- Exec
        if state = x"05" then
          --skip
          state <= x"80";
        else
          if state = x"03" then
            if (ftdcode(31 downto 29) = "001") or (ftdcode(31 downto 30) = "01") or (ftdcode(31 downto 27) = "10001") then
              -- shift,FPU,bf(eq,lt)
              state <= state + 1;
            else
              state <= x"80";
            end if;
          else
            if (state = x"81") and (ftdcode(31 downto 30) < 3) then
              -- without SRAM
              state <= x"FF";
--              state <= x"00";
--              phase <= phase + 1;
            else
              -- with SRAM
              if state = x"8A" then
                --skip
                state <= x"FF";
--                state <= x"00";
--                phase <= phase + 1;
              else
                state <= state + 1;
              end if;
            end if;
          end if;
        end if;
      end if;
      if phase = "100" then
        --skip
        state <= x"00";
        phase <= "000";
--        state <= x"FF";
--        phase <= "111";
      end if;
      if phase = "111" then
        --dummy
        state <= state + 1;
      end if;
      ostate <= "00000000" + state + 1;
    end if;
  end process;
end cocore;

