-- Fetch.vhd
-- Read code from SRAM (Not yet)
-- send back to core.vhd

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity fetch is
  Port (
    clk : in std_logic;
    load_signal : in std_logic := '0';
    pc : in std_logic_vector(31 downto 0);
    inst_sram_request : out std_logic;
    inst_sram_addr : out std_logic_vector(19 downto 0);
    inst_sram_getvalue : in std_logic_vector(31 downto 0);
    inst_sram_request_finished : in std_logic;
    inst_fetched : in std_logic;
    inst : out std_logic_vector(31 downto 0);
    waitwrite : in std_logic_vector(19 downto 0)
  );
end fetch;

architecture fetch_test of fetch is
begin
  fetch_main: process(clk)
  begin
    if rising_edge(clk) then
      if load_signal = '1' then
        if waitwrite = 0 then
if pc = 0 then
	inst <= x"8200F250";
end if;
if pc = 4 then
	inst <= x"43000000";
end if;
if pc = 8 then
	inst <= x"BDCCCCCD";
end if;
if pc = 12 then
	inst <= x"3F666666";
end if;
if pc = 16 then
	inst <= x"3E4CCCCD";
end if;
if pc = 20 then
	inst <= x"C3160000";
end if;
if pc = 24 then
	inst <= x"43160000";
end if;
if pc = 28 then
	inst <= x"3DCCCCCD";
end if;
if pc = 32 then
	inst <= x"C0000000";
end if;
if pc = 36 then
	inst <= x"43800000";
end if;
if pc = 40 then
	inst <= x"4CBEBC20";
end if;
if pc = 44 then
	inst <= x"4E6E6B28";
end if;
if pc = 48 then
	inst <= x"41A00000";
end if;
if pc = 52 then
	inst <= x"3D4CCCCD";
end if;
if pc = 56 then
	inst <= x"3E800000";
end if;
if pc = 60 then
	inst <= x"41200000";
end if;
if pc = 64 then
	inst <= x"3E99999A";
end if;
if pc = 68 then
	inst <= x"437F0000";
end if;
if pc = 72 then
	inst <= x"3E19999A";
end if;
if pc = 76 then
	inst <= x"41700000";
end if;
if pc = 80 then
	inst <= x"40490FDC";
end if;
if pc = 84 then
	inst <= x"41F00000";
end if;
if pc = 88 then
	inst <= x"3C75989E";
end if;
if pc = 92 then
	inst <= x"3F6DA101";
end if;
if pc = 96 then
	inst <= x"3C8F53C5";
end if;
if pc = 100 then
	inst <= x"3E0E9468";
end if;
if pc = 104 then
	inst <= x"3CF30835";
end if;
if pc = 108 then
	inst <= x"38D1B717";
end if;
if pc = 112 then
	inst <= x"BDCCCCCD";
end if;
if pc = 116 then
	inst <= x"3C23D70A";
end if;
if pc = 120 then
	inst <= x"BE4CCCCD";
end if;
if pc = 124 then
	inst <= x"BF800000";
end if;
if pc = 128 then
	inst <= x"40000000";
end if;
if pc = 132 then
	inst <= x"C3480000";
end if;
if pc = 136 then
	inst <= x"43480000";
end if;
if pc = 140 then
	inst <= x"3C8EF998";
end if;
if pc = 144 then
	inst <= x"C0C90FDA";
end if;
if pc = 148 then
	inst <= x"00000000";
end if;
if pc = 152 then
	inst <= x"40C90FDA";
end if;
if pc = 156 then
	inst <= x"3AB39192";
end if;
if pc = 160 then
	inst <= x"3D2AA7DF";
end if;
if pc = 164 then
	inst <= x"3F000000";
end if;
if pc = 168 then
	inst <= x"3F800000";
end if;
if pc = 172 then
	inst <= x"394D8559";
end if;
if pc = 176 then
	inst <= x"3C088723";
end if;
if pc = 180 then
	inst <= x"3E2AAAC1";
end if;
if pc = 184 then
	inst <= x"3F490FD8";
end if;
if pc = 188 then
	inst <= x"3FC90FD8";
end if;
if pc = 192 then
	inst <= x"40490FDC";
end if;
if pc = 196 then
	inst <= x"00000000";
end if;
if pc = 200 then
	inst <= x"00000000";
end if;
if pc = 204 then
	inst <= x"00000000";
end if;
if pc = 208 then
	inst <= x"00000000";
end if;
if pc = 212 then
	inst <= x"00000000";
end if;
if pc = 216 then
	inst <= x"00000000";
end if;
if pc = 220 then
	inst <= x"00000000";
end if;
if pc = 224 then
	inst <= x"00000000";
end if;
if pc = 228 then
	inst <= x"00000000";
end if;
if pc = 232 then
	inst <= x"00000000";
end if;
if pc = 236 then
	inst <= x"00000000";
end if;
if pc = 240 then
	inst <= x"00000000";
end if;
if pc = 244 then
	inst <= x"00000000";
end if;
if pc = 248 then
	inst <= x"00000000";
end if;
if pc = 252 then
	inst <= x"00000000";
end if;
if pc = 256 then
	inst <= x"00000000";
end if;
if pc = 260 then
	inst <= x"00000000";
end if;
if pc = 264 then
	inst <= x"00000000";
end if;
if pc = 268 then
	inst <= x"00000000";
end if;
if pc = 272 then
	inst <= x"00000000";
end if;
if pc = 276 then
	inst <= x"00000000";
end if;
if pc = 280 then
	inst <= x"00000000";
end if;
if pc = 284 then
	inst <= x"00000000";
end if;
if pc = 288 then
	inst <= x"00000000";
end if;
if pc = 292 then
	inst <= x"00000000";
end if;
if pc = 296 then
	inst <= x"00000000";
end if;
if pc = 300 then
	inst <= x"00000000";
end if;
if pc = 304 then
	inst <= x"00000000";
end if;
if pc = 308 then
	inst <= x"00000000";
end if;
if pc = 312 then
	inst <= x"00000000";
end if;
if pc = 316 then
	inst <= x"00000000";
end if;
if pc = 320 then
	inst <= x"00000000";
end if;
if pc = 324 then
	inst <= x"00000000";
end if;
if pc = 328 then
	inst <= x"00000000";
end if;
if pc = 332 then
	inst <= x"00000000";
end if;
if pc = 336 then
	inst <= x"00000000";
end if;
if pc = 340 then
	inst <= x"00000000";
end if;
if pc = 344 then
	inst <= x"00000000";
end if;
if pc = 348 then
	inst <= x"00000000";
end if;
if pc = 352 then
	inst <= x"00000000";
end if;
if pc = 356 then
	inst <= x"00000000";
end if;
if pc = 360 then
	inst <= x"00000000";
end if;
if pc = 364 then
	inst <= x"00000000";
end if;
if pc = 368 then
	inst <= x"00000000";
end if;
if pc = 372 then
	inst <= x"00000000";
end if;
if pc = 376 then
	inst <= x"00000000";
end if;
if pc = 380 then
	inst <= x"00000000";
end if;
if pc = 384 then
	inst <= x"00000000";
end if;
if pc = 388 then
	inst <= x"00000000";
end if;
if pc = 392 then
	inst <= x"00000000";
end if;
if pc = 396 then
	inst <= x"00000000";
end if;
if pc = 400 then
	inst <= x"00000000";
end if;
if pc = 404 then
	inst <= x"00000000";
end if;
if pc = 408 then
	inst <= x"00000000";
end if;
if pc = 412 then
	inst <= x"00000000";
end if;
if pc = 416 then
	inst <= x"00000000";
end if;
if pc = 420 then
	inst <= x"00000000";
end if;
if pc = 424 then
	inst <= x"00000000";
end if;
if pc = 428 then
	inst <= x"00000000";
end if;
if pc = 432 then
	inst <= x"00000000";
end if;
if pc = 436 then
	inst <= x"00000000";
end if;
if pc = 440 then
	inst <= x"00000000";
end if;
if pc = 444 then
	inst <= x"00000000";
end if;
if pc = 448 then
	inst <= x"00000000";
end if;
if pc = 452 then
	inst <= x"00000000";
end if;
if pc = 456 then
	inst <= x"00000000";
end if;
if pc = 460 then
	inst <= x"00000000";
end if;
if pc = 464 then
	inst <= x"00000000";
end if;
if pc = 468 then
	inst <= x"00000000";
end if;
if pc = 472 then
	inst <= x"00000000";
end if;
if pc = 476 then
	inst <= x"437F0000";
end if;
if pc = 480 then
	inst <= x"00000000";
end if;
if pc = 484 then
	inst <= x"00000000";
end if;
if pc = 488 then
	inst <= x"00000000";
end if;
if pc = 492 then
	inst <= x"00000000";
end if;
if pc = 496 then
	inst <= x"00000000";
end if;
if pc = 500 then
	inst <= x"00000000";
end if;
if pc = 504 then
	inst <= x"00000000";
end if;
if pc = 508 then
	inst <= x"00000000";
end if;
if pc = 512 then
	inst <= x"00000000";
end if;
if pc = 516 then
	inst <= x"00000000";
end if;
if pc = 520 then
	inst <= x"00000000";
end if;
if pc = 524 then
	inst <= x"00000000";
end if;
if pc = 528 then
	inst <= x"00000000";
end if;
if pc = 532 then
	inst <= x"00000000";
end if;
if pc = 536 then
	inst <= x"00000000";
end if;
if pc = 540 then
	inst <= x"00000000";
end if;
if pc = 544 then
	inst <= x"00000000";
end if;
if pc = 548 then
	inst <= x"00000000";
end if;
if pc = 552 then
	inst <= x"00000000";
end if;
if pc = 556 then
	inst <= x"00000000";
end if;
if pc = 560 then
	inst <= x"00000000";
end if;
if pc = 564 then
	inst <= x"00000000";
end if;
if pc = 568 then
	inst <= x"00000000";
end if;
if pc = 572 then
	inst <= x"00000000";
end if;
if pc = 576 then
	inst <= x"00000000";
end if;
if pc = 580 then
	inst <= x"00000000";
end if;
if pc = 584 then
	inst <= x"00000000";
end if;
if pc = 588 then
	inst <= x"00000000";
end if;
if pc = 592 then
	inst <= x"00000000";
end if;
if pc = 596 then
	inst <= x"00000000";
end if;
if pc = 600 then
	inst <= x"00000000";
end if;
if pc = 604 then
	inst <= x"00000000";
end if;
if pc = 608 then
	inst <= x"00000000";
end if;
if pc = 612 then
	inst <= x"00000000";
end if;
if pc = 616 then
	inst <= x"00000000";
end if;
if pc = 620 then
	inst <= x"00000000";
end if;
if pc = 624 then
	inst <= x"00000000";
end if;
if pc = 628 then
	inst <= x"00000000";
end if;
if pc = 632 then
	inst <= x"00000000";
end if;
if pc = 636 then
	inst <= x"00000000";
end if;
if pc = 640 then
	inst <= x"00000000";
end if;
if pc = 644 then
	inst <= x"00000000";
end if;
if pc = 648 then
	inst <= x"00000000";
end if;
if pc = 652 then
	inst <= x"00000000";
end if;
if pc = 656 then
	inst <= x"00000000";
end if;
if pc = 660 then
	inst <= x"00000000";
end if;
if pc = 664 then
	inst <= x"00000000";
end if;
if pc = 668 then
	inst <= x"00000000";
end if;
if pc = 672 then
	inst <= x"00000000";
end if;
if pc = 676 then
	inst <= x"00000000";
end if;
if pc = 680 then
	inst <= x"00000000";
end if;
if pc = 684 then
	inst <= x"00000000";
end if;
if pc = 688 then
	inst <= x"00000000";
end if;
if pc = 692 then
	inst <= x"4E6E6B28";
end if;
if pc = 696 then
	inst <= x"00000000";
end if;
if pc = 700 then
	inst <= x"00000000";
end if;
if pc = 704 then
	inst <= x"00000000";
end if;
if pc = 708 then
	inst <= x"00000000";
end if;
if pc = 712 then
	inst <= x"00000000";
end if;
if pc = 716 then
	inst <= x"00000000";
end if;
if pc = 720 then
	inst <= x"00000000";
end if;
if pc = 724 then
	inst <= x"00000000";
end if;
if pc = 728 then
	inst <= x"00000000";
end if;
if pc = 732 then
	inst <= x"00000000";
end if;
if pc = 736 then
	inst <= x"00000000";
end if;
if pc = 740 then
	inst <= x"00000000";
end if;
if pc = 744 then
	inst <= x"00000000";
end if;
if pc = 748 then
	inst <= x"00000000";
end if;
if pc = 752 then
	inst <= x"00000000";
end if;
if pc = 756 then
	inst <= x"00000000";
end if;
if pc = 760 then
	inst <= x"00000000";
end if;
if pc = 764 then
	inst <= x"00000000";
end if;
if pc = 768 then
	inst <= x"00000000";
end if;
if pc = 772 then
	inst <= x"00000000";
end if;
if pc = 776 then
	inst <= x"00000000";
end if;
if pc = 780 then
	inst <= x"00000000";
end if;
if pc = 784 then
	inst <= x"00000000";
end if;
if pc = 788 then
	inst <= x"00000000";
end if;
if pc = 792 then
	inst <= x"00000000";
end if;
if pc = 796 then
	inst <= x"00000000";
end if;
if pc = 800 then
	inst <= x"00000000";
end if;
if pc = 804 then
	inst <= x"00000000";
end if;
if pc = 808 then
	inst <= x"00000000";
end if;
if pc = 812 then
	inst <= x"00000000";
end if;
if pc = 816 then
	inst <= x"00000000";
end if;
if pc = 820 then
	inst <= x"00000000";
end if;
if pc = 824 then
	inst <= x"00000000";
end if;
if pc = 828 then
	inst <= x"00000000";
end if;
if pc = 832 then
	inst <= x"00000000";
end if;
if pc = 836 then
	inst <= x"00000000";
end if;
if pc = 840 then
	inst <= x"00000000";
end if;
if pc = 844 then
	inst <= x"00000000";
end if;
if pc = 848 then
	inst <= x"00000000";
end if;
if pc = 852 then
	inst <= x"00000000";
end if;
if pc = 856 then
	inst <= x"00000000";
end if;
if pc = 860 then
	inst <= x"00000000";
end if;
if pc = 864 then
	inst <= x"00000000";
end if;
if pc = 868 then
	inst <= x"00000000";
end if;
if pc = 872 then
	inst <= x"00000000";
end if;
if pc = 876 then
	inst <= x"00000000";
end if;
if pc = 880 then
	inst <= x"00000000";
end if;
if pc = 884 then
	inst <= x"00000000";
end if;
if pc = 888 then
	inst <= x"00000000";
end if;
if pc = 892 then
	inst <= x"00000000";
end if;
if pc = 896 then
	inst <= x"00000000";
end if;
if pc = 900 then
	inst <= x"00000000";
end if;
if pc = 904 then
	inst <= x"00000000";
end if;
if pc = 908 then
	inst <= x"00000000";
end if;
if pc = 912 then
	inst <= x"00000000";
end if;
if pc = 916 then
	inst <= x"00000000";
end if;
if pc = 920 then
	inst <= x"00000000";
end if;
if pc = 924 then
	inst <= x"00000000";
end if;
if pc = 928 then
	inst <= x"00000000";
end if;
if pc = 932 then
	inst <= x"00000000";
end if;
if pc = 936 then
	inst <= x"00000000";
end if;
if pc = 940 then
	inst <= x"00000000";
end if;
if pc = 944 then
	inst <= x"00000000";
end if;
if pc = 948 then
	inst <= x"00000000";
end if;
if pc = 952 then
	inst <= x"00000000";
end if;
if pc = 956 then
	inst <= x"00000000";
end if;
if pc = 960 then
	inst <= x"00000000";
end if;
if pc = 964 then
	inst <= x"00000000";
end if;
if pc = 968 then
	inst <= x"00000000";
end if;
if pc = 972 then
	inst <= x"00000000";
end if;
if pc = 976 then
	inst <= x"00000000";
end if;
if pc = 980 then
	inst <= x"00000000";
end if;
if pc = 984 then
	inst <= x"00000000";
end if;
if pc = 988 then
	inst <= x"00000000";
end if;
if pc = 992 then
	inst <= x"00000000";
end if;
if pc = 996 then
	inst <= x"00000000";
end if;
if pc = 1000 then
	inst <= x"00000000";
end if;
if pc = 1004 then
	inst <= x"00000000";
end if;
if pc = 1008 then
	inst <= x"00000000";
end if;
if pc = 1012 then
	inst <= x"00000000";
end if;
if pc = 1016 then
	inst <= x"00000000";
end if;
if pc = 1020 then
	inst <= x"00000000";
end if;
if pc = 1024 then
	inst <= x"00000000";
end if;
if pc = 1028 then
	inst <= x"00000000";
end if;
if pc = 1032 then
	inst <= x"00000000";
end if;
if pc = 1036 then
	inst <= x"00000000";
end if;
if pc = 1040 then
	inst <= x"00000000";
end if;
if pc = 1044 then
	inst <= x"00000000";
end if;
if pc = 1048 then
	inst <= x"00000000";
end if;
if pc = 1052 then
	inst <= x"00000000";
end if;
if pc = 1056 then
	inst <= x"00000000";
end if;
if pc = 1060 then
	inst <= x"00000000";
end if;
if pc = 1064 then
	inst <= x"00000000";
end if;
if pc = 1068 then
	inst <= x"00000000";
end if;
if pc = 1072 then
	inst <= x"00000000";
end if;
if pc = 1076 then
	inst <= x"00000000";
end if;
if pc = 1080 then
	inst <= x"00000000";
end if;
if pc = 1084 then
	inst <= x"00000000";
end if;
if pc = 1088 then
	inst <= x"00000000";
end if;
if pc = 1092 then
	inst <= x"00000000";
end if;
if pc = 1096 then
	inst <= x"00000000";
end if;
if pc = 1100 then
	inst <= x"00000000";
end if;
if pc = 1104 then
	inst <= x"00000000";
end if;
if pc = 1108 then
	inst <= x"00000000";
end if;
if pc = 1112 then
	inst <= x"00000000";
end if;
if pc = 1116 then
	inst <= x"00000000";
end if;
if pc = 1120 then
	inst <= x"00000000";
end if;
if pc = 1124 then
	inst <= x"00000000";
end if;
if pc = 1128 then
	inst <= x"00000000";
end if;
if pc = 1132 then
	inst <= x"00000000";
end if;
if pc = 1136 then
	inst <= x"00000000";
end if;
if pc = 1140 then
	inst <= x"00000000";
end if;
if pc = 1144 then
	inst <= x"00000000";
end if;
if pc = 1148 then
	inst <= x"00000000";
end if;
if pc = 1152 then
	inst <= x"00000000";
end if;
if pc = 1156 then
	inst <= x"00000000";
end if;
if pc = 1160 then
	inst <= x"00000000";
end if;
if pc = 1164 then
	inst <= x"00000000";
end if;
if pc = 1168 then
	inst <= x"00000000";
end if;
if pc = 1172 then
	inst <= x"00000000";
end if;
if pc = 1176 then
	inst <= x"00000000";
end if;
if pc = 1180 then
	inst <= x"00000000";
end if;
if pc = 1184 then
	inst <= x"00000000";
end if;
if pc = 1188 then
	inst <= x"00000000";
end if;
if pc = 1192 then
	inst <= x"00000000";
end if;
if pc = 1196 then
	inst <= x"00000000";
end if;
if pc = 1200 then
	inst <= x"00000000";
end if;
if pc = 1204 then
	inst <= x"00000000";
end if;
if pc = 1208 then
	inst <= x"00000000";
end if;
if pc = 1212 then
	inst <= x"00000000";
end if;
if pc = 1216 then
	inst <= x"00000000";
end if;
if pc = 1220 then
	inst <= x"00000000";
end if;
if pc = 1224 then
	inst <= x"00000000";
end if;
if pc = 1228 then
	inst <= x"00000000";
end if;
if pc = 1232 then
	inst <= x"00000000";
end if;
if pc = 1236 then
	inst <= x"00000000";
end if;
if pc = 1240 then
	inst <= x"00000000";
end if;
if pc = 1244 then
	inst <= x"00000000";
end if;
if pc = 1248 then
	inst <= x"00000000";
end if;
if pc = 1252 then
	inst <= x"00000000";
end if;
if pc = 1256 then
	inst <= x"00000000";
end if;
if pc = 1260 then
	inst <= x"00000000";
end if;
if pc = 1264 then
	inst <= x"00000000";
end if;
if pc = 1268 then
	inst <= x"00000000";
end if;
if pc = 1272 then
	inst <= x"00000000";
end if;
if pc = 1276 then
	inst <= x"00000000";
end if;
if pc = 1280 then
	inst <= x"00000000";
end if;
if pc = 1284 then
	inst <= x"00000000";
end if;
if pc = 1288 then
	inst <= x"00000000";
end if;
if pc = 1292 then
	inst <= x"00000000";
end if;
if pc = 1296 then
	inst <= x"00000000";
end if;
if pc = 1300 then
	inst <= x"00000000";
end if;
if pc = 1304 then
	inst <= x"00000000";
end if;
if pc = 1308 then
	inst <= x"00000000";
end if;
if pc = 1312 then
	inst <= x"00000000";
end if;
if pc = 1316 then
	inst <= x"00000000";
end if;
if pc = 1320 then
	inst <= x"00000000";
end if;
if pc = 1324 then
	inst <= x"00000000";
end if;
if pc = 1328 then
	inst <= x"00000000";
end if;
if pc = 1332 then
	inst <= x"00000000";
end if;
if pc = 1336 then
	inst <= x"00000000";
end if;
if pc = 1340 then
	inst <= x"00000000";
end if;
if pc = 1344 then
	inst <= x"00000000";
end if;
if pc = 1348 then
	inst <= x"00000000";
end if;
if pc = 1352 then
	inst <= x"00000000";
end if;
if pc = 1356 then
	inst <= x"00000000";
end if;
if pc = 1360 then
	inst <= x"00000000";
end if;
if pc = 1364 then
	inst <= x"00000000";
end if;
if pc = 1368 then
	inst <= x"00000000";
end if;
if pc = 1372 then
	inst <= x"00000000";
end if;
if pc = 1376 then
	inst <= x"00000000";
end if;
if pc = 1380 then
	inst <= x"00000000";
end if;
if pc = 1384 then
	inst <= x"00000000";
end if;
if pc = 1388 then
	inst <= x"00000000";
end if;
if pc = 1392 then
	inst <= x"00000000";
end if;
if pc = 1396 then
	inst <= x"00000000";
end if;
if pc = 1400 then
	inst <= x"00000000";
end if;
if pc = 1404 then
	inst <= x"00000000";
end if;
if pc = 1408 then
	inst <= x"00000000";
end if;
if pc = 1412 then
	inst <= x"00000000";
end if;
if pc = 1416 then
	inst <= x"00000000";
end if;
if pc = 1420 then
	inst <= x"00000000";
end if;
if pc = 1424 then
	inst <= x"00000000";
end if;
if pc = 1428 then
	inst <= x"00000000";
end if;
if pc = 1432 then
	inst <= x"00000000";
end if;
if pc = 1436 then
	inst <= x"00000000";
end if;
if pc = 1440 then
	inst <= x"00000000";
end if;
if pc = 1444 then
	inst <= x"00000000";
end if;
if pc = 1448 then
	inst <= x"00000000";
end if;
if pc = 1452 then
	inst <= x"00000000";
end if;
if pc = 1456 then
	inst <= x"00000000";
end if;
if pc = 1460 then
	inst <= x"00000000";
end if;
if pc = 1464 then
	inst <= x"00000000";
end if;
if pc = 1468 then
	inst <= x"00000000";
end if;
if pc = 1472 then
	inst <= x"00000000";
end if;
if pc = 1476 then
	inst <= x"00000000";
end if;
if pc = 1480 then
	inst <= x"00000000";
end if;
if pc = 1484 then
	inst <= x"00000000";
end if;
if pc = 1488 then
	inst <= x"00000000";
end if;
if pc = 1492 then
	inst <= x"00000000";
end if;
if pc = 1496 then
	inst <= x"00000000";
end if;
if pc = 1500 then
	inst <= x"00000000";
end if;
if pc = 1504 then
	inst <= x"00000000";
end if;
if pc = 1508 then
	inst <= x"00000000";
end if;
if pc = 1512 then
	inst <= x"00000000";
end if;
if pc = 1516 then
	inst <= x"00000000";
end if;
if pc = 1520 then
	inst <= x"00000000";
end if;
if pc = 1524 then
	inst <= x"00000000";
end if;
if pc = 1528 then
	inst <= x"00000000";
end if;
if pc = 1532 then
	inst <= x"00000000";
end if;
if pc = 1536 then
	inst <= x"00000000";
end if;
if pc = 1540 then
	inst <= x"00000000";
end if;
if pc = 1544 then
	inst <= x"00000000";
end if;
if pc = 1548 then
	inst <= x"00000000";
end if;
if pc = 1552 then
	inst <= x"00000000";
end if;
if pc = 1556 then
	inst <= x"00000000";
end if;
if pc = 1560 then
	inst <= x"00000000";
end if;
if pc = 1564 then
	inst <= x"00000000";
end if;
if pc = 1568 then
	inst <= x"00000000";
end if;
if pc = 1572 then
	inst <= x"00000000";
end if;
if pc = 1576 then
	inst <= x"00000000";
end if;
if pc = 1580 then
	inst <= x"00000000";
end if;
if pc = 1584 then
	inst <= x"00000000";
end if;
if pc = 1588 then
	inst <= x"00000000";
end if;
if pc = 1592 then
	inst <= x"00000000";
end if;
if pc = 1596 then
	inst <= x"00000000";
end if;
if pc = 1600 then
	inst <= x"00000000";
end if;
if pc = 1604 then
	inst <= x"028000EC";
end if;
if pc = 1608 then
	inst <= x"02A000C8";
end if;
if pc = 1612 then
	inst <= x"06C00001";
end if;
if pc = 1616 then
	inst <= x"0220000B";
end if;
if pc = 1620 then
	inst <= x"02400000";
end if;
if pc = 1624 then
	inst <= x"03DC0004";
end if;
if pc = 1628 then
	inst <= x"037E000C";
end if;
if pc = 1632 then
	inst <= x"C57DFFFC";
end if;
if pc = 1636 then
	inst <= x"8200081C";
end if;
if pc = 1640 then
	inst <= x"07DC0004";
end if;
if pc = 1644 then
	inst <= x"0048A000";
end if;
if pc = 1648 then
	inst <= x"C4240000";
end if;
if pc = 1652 then
	inst <= x"06880004";
end if;
if pc = 1656 then
	inst <= x"86C80650";
end if;
if pc = 1660 then
	inst <= x"028000C4";
end if;
if pc = 1664 then
	inst <= x"02A001E0";
end if;
if pc = 1668 then
	inst <= x"02200001";
end if;
if pc = 1672 then
	inst <= x"0240FFFF";
end if;
if pc = 1676 then
	inst <= x"03DC0004";
end if;
if pc = 1680 then
	inst <= x"037E000C";
end if;
if pc = 1684 then
	inst <= x"C57DFFFC";
end if;
if pc = 1688 then
	inst <= x"8200081C";
end if;
if pc = 1692 then
	inst <= x"07DC0004";
end if;
if pc = 1696 then
	inst <= x"0048A000";
end if;
if pc = 1700 then
	inst <= x"C4240000";
end if;
if pc = 1704 then
	inst <= x"06880004";
end if;
if pc = 1708 then
	inst <= x"86C80684";
end if;
if pc = 1712 then
	inst <= x"02200001";
end if;
if pc = 1716 then
	inst <= x"0240FFFF";
end if;
if pc = 1720 then
	inst <= x"03DC0004";
end if;
if pc = 1724 then
	inst <= x"037E000C";
end if;
if pc = 1728 then
	inst <= x"C57DFFFC";
end if;
if pc = 1732 then
	inst <= x"8200081C";
end if;
if pc = 1736 then
	inst <= x"07DC0004";
end if;
if pc = 1740 then
	inst <= x"00420000";
end if;
if pc = 1744 then
	inst <= x"02200001";
end if;
if pc = 1748 then
	inst <= x"03DC0004";
end if;
if pc = 1752 then
	inst <= x"037E000C";
end if;
if pc = 1756 then
	inst <= x"C57DFFFC";
end if;
if pc = 1760 then
	inst <= x"8200081C";
end if;
if pc = 1764 then
	inst <= x"07DC0004";
end if;
if pc = 1768 then
	inst <= x"C42002A8";
end if;
if pc = 1772 then
	inst <= x"02A00368";
end if;
if pc = 1776 then
	inst <= x"02200003";
end if;
if pc = 1780 then
	inst <= x"02400000";
end if;
if pc = 1784 then
	inst <= x"03DC0004";
end if;
if pc = 1788 then
	inst <= x"037E000C";
end if;
if pc = 1792 then
	inst <= x"C57DFFFC";
end if;
if pc = 1796 then
	inst <= x"8200081C";
end if;
if pc = 1800 then
	inst <= x"07DC0004";
end if;
if pc = 1804 then
	inst <= x"C42A0000";
end if;
if pc = 1808 then
	inst <= x"0220003C";
end if;
if pc = 1812 then
	inst <= x"03DC0004";
end if;
if pc = 1816 then
	inst <= x"037E000C";
end if;
if pc = 1820 then
	inst <= x"C57DFFFC";
end if;
if pc = 1824 then
	inst <= x"8200081C";
end if;
if pc = 1828 then
	inst <= x"07DC0004";
end if;
if pc = 1832 then
	inst <= x"C42A0004";
end if;
if pc = 1836 then
	inst <= x"028002CC";
end if;
if pc = 1840 then
	inst <= x"02A00370";
end if;
if pc = 1844 then
	inst <= x"02200002";
end if;
if pc = 1848 then
	inst <= x"03DC0004";
end if;
if pc = 1852 then
	inst <= x"037E000C";
end if;
if pc = 1856 then
	inst <= x"C57DFFFC";
end if;
if pc = 1860 then
	inst <= x"8200081C";
end if;
if pc = 1864 then
	inst <= x"07DC0004";
end if;
if pc = 1868 then
	inst <= x"00E20000";
end if;
if pc = 1872 then
	inst <= x"02200003";
end if;
if pc = 1876 then
	inst <= x"02400000";
end if;
if pc = 1880 then
	inst <= x"03DC0004";
end if;
if pc = 1884 then
	inst <= x"037E000C";
end if;
if pc = 1888 then
	inst <= x"C57DFFFC";
end if;
if pc = 1892 then
	inst <= x"8200081C";
end if;
if pc = 1896 then
	inst <= x"07DC0004";
end if;
if pc = 1900 then
	inst <= x"C4E20004";
end if;
if pc = 1904 then
	inst <= x"0048A000";
end if;
if pc = 1908 then
	inst <= x"C4240000";
end if;
if pc = 1912 then
	inst <= x"06880004";
end if;
if pc = 1916 then
	inst <= x"86C80734";
end if;
if pc = 1920 then
	inst <= x"C1FDFFFC";
end if;
if pc = 1924 then
	inst <= x"E0200000";
end if;
if pc = 1928 then
	inst <= x"C1FDFFFC";
end if;
if pc = 1932 then
	inst <= x"E2200000";
end if;
if pc = 1936 then
	inst <= x"C1FDFFFC";
end if;
if pc = 1940 then
	inst <= x"E0200000";
end if;
if pc = 1944 then
	inst <= x"E0400000";
end if;
if pc = 1948 then
	inst <= x"E0600000";
end if;
if pc = 1952 then
	inst <= x"E0800000";
end if;
if pc = 1956 then
	inst <= x"22221820";
end if;
if pc = 1960 then
	inst <= x"22441020";
end if;
if pc = 1964 then
	inst <= x"22660820";
end if;
if pc = 1968 then
	inst <= x"00224000";
end if;
if pc = 1972 then
	inst <= x"00226000";
end if;
if pc = 1976 then
	inst <= x"00228000";
end if;
if pc = 1980 then
	inst <= x"C1FDFFFC";
end if;
if pc = 1984 then
	inst <= x"E0200000";
end if;
if pc = 1988 then
	inst <= x"E0400000";
end if;
if pc = 1992 then
	inst <= x"E0600000";
end if;
if pc = 1996 then
	inst <= x"E0800000";
end if;
if pc = 2000 then
	inst <= x"22221820";
end if;
if pc = 2004 then
	inst <= x"22441020";
end if;
if pc = 2008 then
	inst <= x"22660820";
end if;
if pc = 2012 then
	inst <= x"00224000";
end if;
if pc = 2016 then
	inst <= x"00226000";
end if;
if pc = 2020 then
	inst <= x"00228000";
end if;
if pc = 2024 then
	inst <= x"C43C0004";
end if;
if pc = 2028 then
	inst <= x"C83C0004";
end if;
if pc = 2032 then
	inst <= x"C1FDFFFC";
end if;
if pc = 2036 then
	inst <= x"CC3C0004";
end if;
if pc = 2040 then
	inst <= x"C03C0004";
end if;
if pc = 2044 then
	inst <= x"228218A0";
end if;
if pc = 2048 then
	inst <= x"226210A0";
end if;
if pc = 2052 then
	inst <= x"224208A0";
end if;
if pc = 2056 then
	inst <= x"E2800000";
end if;
if pc = 2060 then
	inst <= x"E2600000";
end if;
if pc = 2064 then
	inst <= x"E2400000";
end if;
if pc = 2068 then
	inst <= x"E2200000";
end if;
if pc = 2072 then
	inst <= x"C1FDFFFC";
end if;
if pc = 2076 then
	inst <= x"007A0000";
end if;
if pc = 2080 then
	inst <= x"82200834";
end if;
if pc = 2084 then
	inst <= x"C45A0000";
end if;
if pc = 2088 then
	inst <= x"06220001";
end if;
if pc = 2092 then
	inst <= x"03BA0004";
end if;
if pc = 2096 then
	inst <= x"82000820";
end if;
if pc = 2100 then
	inst <= x"00260000";
end if;
if pc = 2104 then
	inst <= x"C1FDFFFC";
end if;
if pc = 2108 then
	inst <= x"50220000";
end if;
if pc = 2112 then
	inst <= x"C1FDFFFC";
end if;
if pc = 2116 then
	inst <= x"60220000";
end if;
if pc = 2120 then
	inst <= x"C1FDFFFC";
end if;
if pc = 2124 then
	inst <= x"C84000C0";
end if;
if pc = 2128 then
	inst <= x"C86000BC";
end if;
if pc = 2132 then
	inst <= x"C88000B8";
end if;
if pc = 2136 then
	inst <= x"C43C0000";
end if;
if pc = 2140 then
	inst <= x"8E240A10";
end if;
if pc = 2144 then
	inst <= x"44224000";
end if;
if pc = 2148 then
	inst <= x"04402000";
end if;
if pc = 2152 then
	inst <= x"C45C0004";
end if;
if pc = 2156 then
	inst <= x"8E240898";
end if;
if pc = 2160 then
	inst <= x"44224000";
end if;
if pc = 2164 then
	inst <= x"04604000";
end if;
if pc = 2168 then
	inst <= x"C17DFFFC";
end if;
if pc = 2172 then
	inst <= x"00260000";
end if;
if pc = 2176 then
	inst <= x"03DC0010";
end if;
if pc = 2180 then
	inst <= x"037E000C";
end if;
if pc = 2184 then
	inst <= x"C57DFFFC";
end if;
if pc = 2188 then
	inst <= x"8200084C";
end if;
if pc = 2192 then
	inst <= x"07DC0010";
end if;
if pc = 2196 then
	inst <= x"820009F8";
end if;
if pc = 2200 then
	inst <= x"8E26094C";
end if;
if pc = 2204 then
	inst <= x"8E8208F8";
end if;
if pc = 2208 then
	inst <= x"C84000B4";
end if;
if pc = 2212 then
	inst <= x"48442000";
end if;
if pc = 2216 then
	inst <= x"48442000";
end if;
if pc = 2220 then
	inst <= x"48442000";
end if;
if pc = 2224 then
	inst <= x"44424000";
end if;
if pc = 2228 then
	inst <= x"C86000B0";
end if;
if pc = 2232 then
	inst <= x"48662000";
end if;
if pc = 2236 then
	inst <= x"48662000";
end if;
if pc = 2240 then
	inst <= x"48662000";
end if;
if pc = 2244 then
	inst <= x"48662000";
end if;
if pc = 2248 then
	inst <= x"48662000";
end if;
if pc = 2252 then
	inst <= x"40446000";
end if;
if pc = 2256 then
	inst <= x"C86000AC";
end if;
if pc = 2260 then
	inst <= x"48662000";
end if;
if pc = 2264 then
	inst <= x"48662000";
end if;
if pc = 2268 then
	inst <= x"48662000";
end if;
if pc = 2272 then
	inst <= x"48662000";
end if;
if pc = 2276 then
	inst <= x"48662000";
end if;
if pc = 2280 then
	inst <= x"48662000";
end if;
if pc = 2284 then
	inst <= x"48262000";
end if;
if pc = 2288 then
	inst <= x"44242000";
end if;
if pc = 2292 then
	inst <= x"82000948";
end if;
if pc = 2296 then
	inst <= x"44262000";
end if;
if pc = 2300 then
	inst <= x"C84000A8";
end if;
if pc = 2304 then
	inst <= x"C86000A4";
end if;
if pc = 2308 then
	inst <= x"48662000";
end if;
if pc = 2312 then
	inst <= x"48662000";
end if;
if pc = 2316 then
	inst <= x"44446000";
end if;
if pc = 2320 then
	inst <= x"C86000A0";
end if;
if pc = 2324 then
	inst <= x"48662000";
end if;
if pc = 2328 then
	inst <= x"48662000";
end if;
if pc = 2332 then
	inst <= x"48662000";
end if;
if pc = 2336 then
	inst <= x"48662000";
end if;
if pc = 2340 then
	inst <= x"40446000";
end if;
if pc = 2344 then
	inst <= x"C860009C";
end if;
if pc = 2348 then
	inst <= x"48662000";
end if;
if pc = 2352 then
	inst <= x"48662000";
end if;
if pc = 2356 then
	inst <= x"48662000";
end if;
if pc = 2360 then
	inst <= x"48662000";
end if;
if pc = 2364 then
	inst <= x"48662000";
end if;
if pc = 2368 then
	inst <= x"48262000";
end if;
if pc = 2372 then
	inst <= x"44242000";
end if;
if pc = 2376 then
	inst <= x"820009F8";
end if;
if pc = 2380 then
	inst <= x"8E8209A8";
end if;
if pc = 2384 then
	inst <= x"C84000B4";
end if;
if pc = 2388 then
	inst <= x"48442000";
end if;
if pc = 2392 then
	inst <= x"48442000";
end if;
if pc = 2396 then
	inst <= x"48442000";
end if;
if pc = 2400 then
	inst <= x"44424000";
end if;
if pc = 2404 then
	inst <= x"C86000B0";
end if;
if pc = 2408 then
	inst <= x"48662000";
end if;
if pc = 2412 then
	inst <= x"48662000";
end if;
if pc = 2416 then
	inst <= x"48662000";
end if;
if pc = 2420 then
	inst <= x"48662000";
end if;
if pc = 2424 then
	inst <= x"48662000";
end if;
if pc = 2428 then
	inst <= x"40446000";
end if;
if pc = 2432 then
	inst <= x"C86000AC";
end if;
if pc = 2436 then
	inst <= x"48662000";
end if;
if pc = 2440 then
	inst <= x"48662000";
end if;
if pc = 2444 then
	inst <= x"48662000";
end if;
if pc = 2448 then
	inst <= x"48662000";
end if;
if pc = 2452 then
	inst <= x"48662000";
end if;
if pc = 2456 then
	inst <= x"48662000";
end if;
if pc = 2460 then
	inst <= x"48262000";
end if;
if pc = 2464 then
	inst <= x"44242000";
end if;
if pc = 2468 then
	inst <= x"820009F8";
end if;
if pc = 2472 then
	inst <= x"44262000";
end if;
if pc = 2476 then
	inst <= x"C84000A8";
end if;
if pc = 2480 then
	inst <= x"C86000A4";
end if;
if pc = 2484 then
	inst <= x"48662000";
end if;
if pc = 2488 then
	inst <= x"48662000";
end if;
if pc = 2492 then
	inst <= x"44446000";
end if;
if pc = 2496 then
	inst <= x"C86000A0";
end if;
if pc = 2500 then
	inst <= x"48662000";
end if;
if pc = 2504 then
	inst <= x"48662000";
end if;
if pc = 2508 then
	inst <= x"48662000";
end if;
if pc = 2512 then
	inst <= x"48662000";
end if;
if pc = 2516 then
	inst <= x"40446000";
end if;
if pc = 2520 then
	inst <= x"C860009C";
end if;
if pc = 2524 then
	inst <= x"48662000";
end if;
if pc = 2528 then
	inst <= x"48662000";
end if;
if pc = 2532 then
	inst <= x"48662000";
end if;
if pc = 2536 then
	inst <= x"48662000";
end if;
if pc = 2540 then
	inst <= x"48662000";
end if;
if pc = 2544 then
	inst <= x"48262000";
end if;
if pc = 2548 then
	inst <= x"44242000";
end if;
if pc = 2552 then
	inst <= x"02200001";
end if;
if pc = 2556 then
	inst <= x"C05C0004";
end if;
if pc = 2560 then
	inst <= x"82420A08";
end if;
if pc = 2564 then
	inst <= x"82000A0C";
end if;
if pc = 2568 then
	inst <= x"44202000";
end if;
if pc = 2572 then
	inst <= x"82000B70";
end if;
if pc = 2576 then
	inst <= x"8E260AC4";
end if;
if pc = 2580 then
	inst <= x"8E820A70";
end if;
if pc = 2584 then
	inst <= x"C84000B4";
end if;
if pc = 2588 then
	inst <= x"48442000";
end if;
if pc = 2592 then
	inst <= x"48442000";
end if;
if pc = 2596 then
	inst <= x"48442000";
end if;
if pc = 2600 then
	inst <= x"44424000";
end if;
if pc = 2604 then
	inst <= x"C86000B0";
end if;
if pc = 2608 then
	inst <= x"48662000";
end if;
if pc = 2612 then
	inst <= x"48662000";
end if;
if pc = 2616 then
	inst <= x"48662000";
end if;
if pc = 2620 then
	inst <= x"48662000";
end if;
if pc = 2624 then
	inst <= x"48662000";
end if;
if pc = 2628 then
	inst <= x"40446000";
end if;
if pc = 2632 then
	inst <= x"C86000AC";
end if;
if pc = 2636 then
	inst <= x"48662000";
end if;
if pc = 2640 then
	inst <= x"48662000";
end if;
if pc = 2644 then
	inst <= x"48662000";
end if;
if pc = 2648 then
	inst <= x"48662000";
end if;
if pc = 2652 then
	inst <= x"48662000";
end if;
if pc = 2656 then
	inst <= x"48662000";
end if;
if pc = 2660 then
	inst <= x"48262000";
end if;
if pc = 2664 then
	inst <= x"44242000";
end if;
if pc = 2668 then
	inst <= x"82000AC0";
end if;
if pc = 2672 then
	inst <= x"44262000";
end if;
if pc = 2676 then
	inst <= x"C84000A8";
end if;
if pc = 2680 then
	inst <= x"C86000A4";
end if;
if pc = 2684 then
	inst <= x"48662000";
end if;
if pc = 2688 then
	inst <= x"48662000";
end if;
if pc = 2692 then
	inst <= x"44446000";
end if;
if pc = 2696 then
	inst <= x"C86000A0";
end if;
if pc = 2700 then
	inst <= x"48662000";
end if;
if pc = 2704 then
	inst <= x"48662000";
end if;
if pc = 2708 then
	inst <= x"48662000";
end if;
if pc = 2712 then
	inst <= x"48662000";
end if;
if pc = 2716 then
	inst <= x"40446000";
end if;
if pc = 2720 then
	inst <= x"C860009C";
end if;
if pc = 2724 then
	inst <= x"48662000";
end if;
if pc = 2728 then
	inst <= x"48662000";
end if;
if pc = 2732 then
	inst <= x"48662000";
end if;
if pc = 2736 then
	inst <= x"48662000";
end if;
if pc = 2740 then
	inst <= x"48662000";
end if;
if pc = 2744 then
	inst <= x"48262000";
end if;
if pc = 2748 then
	inst <= x"44242000";
end if;
if pc = 2752 then
	inst <= x"82000B70";
end if;
if pc = 2756 then
	inst <= x"8E820B20";
end if;
if pc = 2760 then
	inst <= x"C84000B4";
end if;
if pc = 2764 then
	inst <= x"48442000";
end if;
if pc = 2768 then
	inst <= x"48442000";
end if;
if pc = 2772 then
	inst <= x"48442000";
end if;
if pc = 2776 then
	inst <= x"44424000";
end if;
if pc = 2780 then
	inst <= x"C86000B0";
end if;
if pc = 2784 then
	inst <= x"48662000";
end if;
if pc = 2788 then
	inst <= x"48662000";
end if;
if pc = 2792 then
	inst <= x"48662000";
end if;
if pc = 2796 then
	inst <= x"48662000";
end if;
if pc = 2800 then
	inst <= x"48662000";
end if;
if pc = 2804 then
	inst <= x"40446000";
end if;
if pc = 2808 then
	inst <= x"C86000AC";
end if;
if pc = 2812 then
	inst <= x"48662000";
end if;
if pc = 2816 then
	inst <= x"48662000";
end if;
if pc = 2820 then
	inst <= x"48662000";
end if;
if pc = 2824 then
	inst <= x"48662000";
end if;
if pc = 2828 then
	inst <= x"48662000";
end if;
if pc = 2832 then
	inst <= x"48662000";
end if;
if pc = 2836 then
	inst <= x"48262000";
end if;
if pc = 2840 then
	inst <= x"44242000";
end if;
if pc = 2844 then
	inst <= x"82000B70";
end if;
if pc = 2848 then
	inst <= x"44262000";
end if;
if pc = 2852 then
	inst <= x"C84000A8";
end if;
if pc = 2856 then
	inst <= x"C86000A4";
end if;
if pc = 2860 then
	inst <= x"48662000";
end if;
if pc = 2864 then
	inst <= x"48662000";
end if;
if pc = 2868 then
	inst <= x"44446000";
end if;
if pc = 2872 then
	inst <= x"C86000A0";
end if;
if pc = 2876 then
	inst <= x"48662000";
end if;
if pc = 2880 then
	inst <= x"48662000";
end if;
if pc = 2884 then
	inst <= x"48662000";
end if;
if pc = 2888 then
	inst <= x"48662000";
end if;
if pc = 2892 then
	inst <= x"40446000";
end if;
if pc = 2896 then
	inst <= x"C860009C";
end if;
if pc = 2900 then
	inst <= x"48662000";
end if;
if pc = 2904 then
	inst <= x"48662000";
end if;
if pc = 2908 then
	inst <= x"48662000";
end if;
if pc = 2912 then
	inst <= x"48662000";
end if;
if pc = 2916 then
	inst <= x"48662000";
end if;
if pc = 2920 then
	inst <= x"48262000";
end if;
if pc = 2924 then
	inst <= x"44242000";
end if;
if pc = 2928 then
	inst <= x"02200001";
end if;
if pc = 2932 then
	inst <= x"C05C0000";
end if;
if pc = 2936 then
	inst <= x"82420B80";
end if;
if pc = 2940 then
	inst <= x"C1FDFFFC";
end if;
if pc = 2944 then
	inst <= x"44202000";
end if;
if pc = 2948 then
	inst <= x"C1FDFFFC";
end if;
if pc = 2952 then
	inst <= x"C84000C0";
end if;
if pc = 2956 then
	inst <= x"C86000BC";
end if;
if pc = 2960 then
	inst <= x"C88000B8";
end if;
if pc = 2964 then
	inst <= x"C43C0000";
end if;
if pc = 2968 then
	inst <= x"8E240D4C";
end if;
if pc = 2972 then
	inst <= x"44224000";
end if;
if pc = 2976 then
	inst <= x"04402000";
end if;
if pc = 2980 then
	inst <= x"C45C0004";
end if;
if pc = 2984 then
	inst <= x"8E240BD4";
end if;
if pc = 2988 then
	inst <= x"44224000";
end if;
if pc = 2992 then
	inst <= x"04604000";
end if;
if pc = 2996 then
	inst <= x"C17DFFFC";
end if;
if pc = 3000 then
	inst <= x"00260000";
end if;
if pc = 3004 then
	inst <= x"03DC0010";
end if;
if pc = 3008 then
	inst <= x"037E000C";
end if;
if pc = 3012 then
	inst <= x"C57DFFFC";
end if;
if pc = 3016 then
	inst <= x"8200084C";
end if;
if pc = 3020 then
	inst <= x"07DC0010";
end if;
if pc = 3024 then
	inst <= x"82000D34";
end if;
if pc = 3028 then
	inst <= x"8E260C88";
end if;
if pc = 3032 then
	inst <= x"8E820C34";
end if;
if pc = 3036 then
	inst <= x"C84000B4";
end if;
if pc = 3040 then
	inst <= x"48442000";
end if;
if pc = 3044 then
	inst <= x"48442000";
end if;
if pc = 3048 then
	inst <= x"48442000";
end if;
if pc = 3052 then
	inst <= x"44424000";
end if;
if pc = 3056 then
	inst <= x"C86000B0";
end if;
if pc = 3060 then
	inst <= x"48662000";
end if;
if pc = 3064 then
	inst <= x"48662000";
end if;
if pc = 3068 then
	inst <= x"48662000";
end if;
if pc = 3072 then
	inst <= x"48662000";
end if;
if pc = 3076 then
	inst <= x"48662000";
end if;
if pc = 3080 then
	inst <= x"40446000";
end if;
if pc = 3084 then
	inst <= x"C86000AC";
end if;
if pc = 3088 then
	inst <= x"48662000";
end if;
if pc = 3092 then
	inst <= x"48662000";
end if;
if pc = 3096 then
	inst <= x"48662000";
end if;
if pc = 3100 then
	inst <= x"48662000";
end if;
if pc = 3104 then
	inst <= x"48662000";
end if;
if pc = 3108 then
	inst <= x"48662000";
end if;
if pc = 3112 then
	inst <= x"48262000";
end if;
if pc = 3116 then
	inst <= x"44242000";
end if;
if pc = 3120 then
	inst <= x"82000C84";
end if;
if pc = 3124 then
	inst <= x"44262000";
end if;
if pc = 3128 then
	inst <= x"C84000A8";
end if;
if pc = 3132 then
	inst <= x"C86000A4";
end if;
if pc = 3136 then
	inst <= x"48662000";
end if;
if pc = 3140 then
	inst <= x"48662000";
end if;
if pc = 3144 then
	inst <= x"44446000";
end if;
if pc = 3148 then
	inst <= x"C86000A0";
end if;
if pc = 3152 then
	inst <= x"48662000";
end if;
if pc = 3156 then
	inst <= x"48662000";
end if;
if pc = 3160 then
	inst <= x"48662000";
end if;
if pc = 3164 then
	inst <= x"48662000";
end if;
if pc = 3168 then
	inst <= x"40446000";
end if;
if pc = 3172 then
	inst <= x"C860009C";
end if;
if pc = 3176 then
	inst <= x"48662000";
end if;
if pc = 3180 then
	inst <= x"48662000";
end if;
if pc = 3184 then
	inst <= x"48662000";
end if;
if pc = 3188 then
	inst <= x"48662000";
end if;
if pc = 3192 then
	inst <= x"48662000";
end if;
if pc = 3196 then
	inst <= x"48262000";
end if;
if pc = 3200 then
	inst <= x"44242000";
end if;
if pc = 3204 then
	inst <= x"82000D34";
end if;
if pc = 3208 then
	inst <= x"8E820CE4";
end if;
if pc = 3212 then
	inst <= x"C84000B4";
end if;
if pc = 3216 then
	inst <= x"48442000";
end if;
if pc = 3220 then
	inst <= x"48442000";
end if;
if pc = 3224 then
	inst <= x"48442000";
end if;
if pc = 3228 then
	inst <= x"44424000";
end if;
if pc = 3232 then
	inst <= x"C86000B0";
end if;
if pc = 3236 then
	inst <= x"48662000";
end if;
if pc = 3240 then
	inst <= x"48662000";
end if;
if pc = 3244 then
	inst <= x"48662000";
end if;
if pc = 3248 then
	inst <= x"48662000";
end if;
if pc = 3252 then
	inst <= x"48662000";
end if;
if pc = 3256 then
	inst <= x"40446000";
end if;
if pc = 3260 then
	inst <= x"C86000AC";
end if;
if pc = 3264 then
	inst <= x"48662000";
end if;
if pc = 3268 then
	inst <= x"48662000";
end if;
if pc = 3272 then
	inst <= x"48662000";
end if;
if pc = 3276 then
	inst <= x"48662000";
end if;
if pc = 3280 then
	inst <= x"48662000";
end if;
if pc = 3284 then
	inst <= x"48662000";
end if;
if pc = 3288 then
	inst <= x"48262000";
end if;
if pc = 3292 then
	inst <= x"44242000";
end if;
if pc = 3296 then
	inst <= x"82000D34";
end if;
if pc = 3300 then
	inst <= x"44262000";
end if;
if pc = 3304 then
	inst <= x"C84000A8";
end if;
if pc = 3308 then
	inst <= x"C86000A4";
end if;
if pc = 3312 then
	inst <= x"48662000";
end if;
if pc = 3316 then
	inst <= x"48662000";
end if;
if pc = 3320 then
	inst <= x"44446000";
end if;
if pc = 3324 then
	inst <= x"C86000A0";
end if;
if pc = 3328 then
	inst <= x"48662000";
end if;
if pc = 3332 then
	inst <= x"48662000";
end if;
if pc = 3336 then
	inst <= x"48662000";
end if;
if pc = 3340 then
	inst <= x"48662000";
end if;
if pc = 3344 then
	inst <= x"40446000";
end if;
if pc = 3348 then
	inst <= x"C860009C";
end if;
if pc = 3352 then
	inst <= x"48662000";
end if;
if pc = 3356 then
	inst <= x"48662000";
end if;
if pc = 3360 then
	inst <= x"48662000";
end if;
if pc = 3364 then
	inst <= x"48662000";
end if;
if pc = 3368 then
	inst <= x"48662000";
end if;
if pc = 3372 then
	inst <= x"48262000";
end if;
if pc = 3376 then
	inst <= x"44242000";
end if;
if pc = 3380 then
	inst <= x"02200001";
end if;
if pc = 3384 then
	inst <= x"C05C0004";
end if;
if pc = 3388 then
	inst <= x"82420D44";
end if;
if pc = 3392 then
	inst <= x"82000D48";
end if;
if pc = 3396 then
	inst <= x"44202000";
end if;
if pc = 3400 then
	inst <= x"82000EAC";
end if;
if pc = 3404 then
	inst <= x"8E260E00";
end if;
if pc = 3408 then
	inst <= x"8E820DA4";
end if;
if pc = 3412 then
	inst <= x"C84000A8";
end if;
if pc = 3416 then
	inst <= x"C86000A4";
end if;
if pc = 3420 then
	inst <= x"48662000";
end if;
if pc = 3424 then
	inst <= x"48662000";
end if;
if pc = 3428 then
	inst <= x"44446000";
end if;
if pc = 3432 then
	inst <= x"C86000A0";
end if;
if pc = 3436 then
	inst <= x"48662000";
end if;
if pc = 3440 then
	inst <= x"48662000";
end if;
if pc = 3444 then
	inst <= x"48662000";
end if;
if pc = 3448 then
	inst <= x"48662000";
end if;
if pc = 3452 then
	inst <= x"40446000";
end if;
if pc = 3456 then
	inst <= x"C860009C";
end if;
if pc = 3460 then
	inst <= x"48662000";
end if;
if pc = 3464 then
	inst <= x"48662000";
end if;
if pc = 3468 then
	inst <= x"48662000";
end if;
if pc = 3472 then
	inst <= x"48662000";
end if;
if pc = 3476 then
	inst <= x"48662000";
end if;
if pc = 3480 then
	inst <= x"48262000";
end if;
if pc = 3484 then
	inst <= x"44242000";
end if;
if pc = 3488 then
	inst <= x"82000DFC";
end if;
if pc = 3492 then
	inst <= x"44262000";
end if;
if pc = 3496 then
	inst <= x"C84000B4";
end if;
if pc = 3500 then
	inst <= x"48442000";
end if;
if pc = 3504 then
	inst <= x"48442000";
end if;
if pc = 3508 then
	inst <= x"48442000";
end if;
if pc = 3512 then
	inst <= x"44424000";
end if;
if pc = 3516 then
	inst <= x"C86000B0";
end if;
if pc = 3520 then
	inst <= x"48662000";
end if;
if pc = 3524 then
	inst <= x"48662000";
end if;
if pc = 3528 then
	inst <= x"48662000";
end if;
if pc = 3532 then
	inst <= x"48662000";
end if;
if pc = 3536 then
	inst <= x"48662000";
end if;
if pc = 3540 then
	inst <= x"40446000";
end if;
if pc = 3544 then
	inst <= x"C86000AC";
end if;
if pc = 3548 then
	inst <= x"48662000";
end if;
if pc = 3552 then
	inst <= x"48662000";
end if;
if pc = 3556 then
	inst <= x"48662000";
end if;
if pc = 3560 then
	inst <= x"48662000";
end if;
if pc = 3564 then
	inst <= x"48662000";
end if;
if pc = 3568 then
	inst <= x"48662000";
end if;
if pc = 3572 then
	inst <= x"48262000";
end if;
if pc = 3576 then
	inst <= x"44242000";
end if;
if pc = 3580 then
	inst <= x"82000EAC";
end if;
if pc = 3584 then
	inst <= x"8E820E54";
end if;
if pc = 3588 then
	inst <= x"C84000A8";
end if;
if pc = 3592 then
	inst <= x"C86000A4";
end if;
if pc = 3596 then
	inst <= x"48662000";
end if;
if pc = 3600 then
	inst <= x"48662000";
end if;
if pc = 3604 then
	inst <= x"44446000";
end if;
if pc = 3608 then
	inst <= x"C86000A0";
end if;
if pc = 3612 then
	inst <= x"48662000";
end if;
if pc = 3616 then
	inst <= x"48662000";
end if;
if pc = 3620 then
	inst <= x"48662000";
end if;
if pc = 3624 then
	inst <= x"48662000";
end if;
if pc = 3628 then
	inst <= x"40446000";
end if;
if pc = 3632 then
	inst <= x"C860009C";
end if;
if pc = 3636 then
	inst <= x"48662000";
end if;
if pc = 3640 then
	inst <= x"48662000";
end if;
if pc = 3644 then
	inst <= x"48662000";
end if;
if pc = 3648 then
	inst <= x"48662000";
end if;
if pc = 3652 then
	inst <= x"48662000";
end if;
if pc = 3656 then
	inst <= x"48262000";
end if;
if pc = 3660 then
	inst <= x"44242000";
end if;
if pc = 3664 then
	inst <= x"82000EAC";
end if;
if pc = 3668 then
	inst <= x"44262000";
end if;
if pc = 3672 then
	inst <= x"C84000B4";
end if;
if pc = 3676 then
	inst <= x"48442000";
end if;
if pc = 3680 then
	inst <= x"48442000";
end if;
if pc = 3684 then
	inst <= x"48442000";
end if;
if pc = 3688 then
	inst <= x"44424000";
end if;
if pc = 3692 then
	inst <= x"C86000B0";
end if;
if pc = 3696 then
	inst <= x"48662000";
end if;
if pc = 3700 then
	inst <= x"48662000";
end if;
if pc = 3704 then
	inst <= x"48662000";
end if;
if pc = 3708 then
	inst <= x"48662000";
end if;
if pc = 3712 then
	inst <= x"48662000";
end if;
if pc = 3716 then
	inst <= x"40446000";
end if;
if pc = 3720 then
	inst <= x"C86000AC";
end if;
if pc = 3724 then
	inst <= x"48662000";
end if;
if pc = 3728 then
	inst <= x"48662000";
end if;
if pc = 3732 then
	inst <= x"48662000";
end if;
if pc = 3736 then
	inst <= x"48662000";
end if;
if pc = 3740 then
	inst <= x"48662000";
end if;
if pc = 3744 then
	inst <= x"48662000";
end if;
if pc = 3748 then
	inst <= x"48262000";
end if;
if pc = 3752 then
	inst <= x"44242000";
end if;
if pc = 3756 then
	inst <= x"02200001";
end if;
if pc = 3760 then
	inst <= x"C05C0000";
end if;
if pc = 3764 then
	inst <= x"82420EBC";
end if;
if pc = 3768 then
	inst <= x"C1FDFFFC";
end if;
if pc = 3772 then
	inst <= x"44202000";
end if;
if pc = 3776 then
	inst <= x"C1FDFFFC";
end if;
if pc = 3780 then
	inst <= x"C8400098";
end if;
if pc = 3784 then
	inst <= x"8E240F00";
end if;
if pc = 3788 then
	inst <= x"44224000";
end if;
if pc = 3792 then
	inst <= x"8E240EDC";
end if;
if pc = 3796 then
	inst <= x"44224000";
end if;
if pc = 3800 then
	inst <= x"82000EC4";
end if;
if pc = 3804 then
	inst <= x"8E020EF8";
end if;
if pc = 3808 then
	inst <= x"C8600090";
end if;
if pc = 3812 then
	inst <= x"8E620EF0";
end if;
if pc = 3816 then
	inst <= x"40224000";
end if;
if pc = 3820 then
	inst <= x"82000EC4";
end if;
if pc = 3824 then
	inst <= x"02200001";
end if;
if pc = 3828 then
	inst <= x"8200084C";
end if;
if pc = 3832 then
	inst <= x"0220FFFF";
end if;
if pc = 3836 then
	inst <= x"8200084C";
end if;
if pc = 3840 then
	inst <= x"8E0210D8";
end if;
if pc = 3844 then
	inst <= x"C8600090";
end if;
if pc = 3848 then
	inst <= x"8E620F3C";
end if;
if pc = 3852 then
	inst <= x"40224000";
end if;
if pc = 3856 then
	inst <= x"8E240F1C";
end if;
if pc = 3860 then
	inst <= x"44224000";
end if;
if pc = 3864 then
	inst <= x"82000EC4";
end if;
if pc = 3868 then
	inst <= x"8E020F34";
end if;
if pc = 3872 then
	inst <= x"8E620F2C";
end if;
if pc = 3876 then
	inst <= x"40224000";
end if;
if pc = 3880 then
	inst <= x"82000EC4";
end if;
if pc = 3884 then
	inst <= x"02200001";
end if;
if pc = 3888 then
	inst <= x"8200084C";
end if;
if pc = 3892 then
	inst <= x"0220FFFF";
end if;
if pc = 3896 then
	inst <= x"8200084C";
end if;
if pc = 3900 then
	inst <= x"C84000C0";
end if;
if pc = 3904 then
	inst <= x"C86000BC";
end if;
if pc = 3908 then
	inst <= x"C88000B8";
end if;
if pc = 3912 then
	inst <= x"8E240F70";
end if;
if pc = 3916 then
	inst <= x"44224000";
end if;
if pc = 3920 then
	inst <= x"0220FFFF";
end if;
if pc = 3924 then
	inst <= x"C17DFFFC";
end if;
if pc = 3928 then
	inst <= x"03DC0008";
end if;
if pc = 3932 then
	inst <= x"037E000C";
end if;
if pc = 3936 then
	inst <= x"C57DFFFC";
end if;
if pc = 3940 then
	inst <= x"8200084C";
end if;
if pc = 3944 then
	inst <= x"07DC0008";
end if;
if pc = 3948 then
	inst <= x"820010D0";
end if;
if pc = 3952 then
	inst <= x"8E261024";
end if;
if pc = 3956 then
	inst <= x"8E820FD0";
end if;
if pc = 3960 then
	inst <= x"C84000B4";
end if;
if pc = 3964 then
	inst <= x"48442000";
end if;
if pc = 3968 then
	inst <= x"48442000";
end if;
if pc = 3972 then
	inst <= x"48442000";
end if;
if pc = 3976 then
	inst <= x"44424000";
end if;
if pc = 3980 then
	inst <= x"C86000B0";
end if;
if pc = 3984 then
	inst <= x"48662000";
end if;
if pc = 3988 then
	inst <= x"48662000";
end if;
if pc = 3992 then
	inst <= x"48662000";
end if;
if pc = 3996 then
	inst <= x"48662000";
end if;
if pc = 4000 then
	inst <= x"48662000";
end if;
if pc = 4004 then
	inst <= x"40446000";
end if;
if pc = 4008 then
	inst <= x"C86000AC";
end if;
if pc = 4012 then
	inst <= x"48662000";
end if;
if pc = 4016 then
	inst <= x"48662000";
end if;
if pc = 4020 then
	inst <= x"48662000";
end if;
if pc = 4024 then
	inst <= x"48662000";
end if;
if pc = 4028 then
	inst <= x"48662000";
end if;
if pc = 4032 then
	inst <= x"48662000";
end if;
if pc = 4036 then
	inst <= x"48262000";
end if;
if pc = 4040 then
	inst <= x"44242000";
end if;
if pc = 4044 then
	inst <= x"82001020";
end if;
if pc = 4048 then
	inst <= x"44262000";
end if;
if pc = 4052 then
	inst <= x"C84000A8";
end if;
if pc = 4056 then
	inst <= x"C86000A4";
end if;
if pc = 4060 then
	inst <= x"48662000";
end if;
if pc = 4064 then
	inst <= x"48662000";
end if;
if pc = 4068 then
	inst <= x"44446000";
end if;
if pc = 4072 then
	inst <= x"C86000A0";
end if;
if pc = 4076 then
	inst <= x"48662000";
end if;
if pc = 4080 then
	inst <= x"48662000";
end if;
if pc = 4084 then
	inst <= x"48662000";
end if;
if pc = 4088 then
	inst <= x"48662000";
end if;
if pc = 4092 then
	inst <= x"40446000";
end if;
if pc = 4096 then
	inst <= x"C860009C";
end if;
if pc = 4100 then
	inst <= x"48662000";
end if;
if pc = 4104 then
	inst <= x"48662000";
end if;
if pc = 4108 then
	inst <= x"48662000";
end if;
if pc = 4112 then
	inst <= x"48662000";
end if;
if pc = 4116 then
	inst <= x"48662000";
end if;
if pc = 4120 then
	inst <= x"48262000";
end if;
if pc = 4124 then
	inst <= x"44242000";
end if;
if pc = 4128 then
	inst <= x"820010D0";
end if;
if pc = 4132 then
	inst <= x"8E821080";
end if;
if pc = 4136 then
	inst <= x"C84000B4";
end if;
if pc = 4140 then
	inst <= x"48442000";
end if;
if pc = 4144 then
	inst <= x"48442000";
end if;
if pc = 4148 then
	inst <= x"48442000";
end if;
if pc = 4152 then
	inst <= x"44424000";
end if;
if pc = 4156 then
	inst <= x"C86000B0";
end if;
if pc = 4160 then
	inst <= x"48662000";
end if;
if pc = 4164 then
	inst <= x"48662000";
end if;
if pc = 4168 then
	inst <= x"48662000";
end if;
if pc = 4172 then
	inst <= x"48662000";
end if;
if pc = 4176 then
	inst <= x"48662000";
end if;
if pc = 4180 then
	inst <= x"40446000";
end if;
if pc = 4184 then
	inst <= x"C86000AC";
end if;
if pc = 4188 then
	inst <= x"48662000";
end if;
if pc = 4192 then
	inst <= x"48662000";
end if;
if pc = 4196 then
	inst <= x"48662000";
end if;
if pc = 4200 then
	inst <= x"48662000";
end if;
if pc = 4204 then
	inst <= x"48662000";
end if;
if pc = 4208 then
	inst <= x"48662000";
end if;
if pc = 4212 then
	inst <= x"48262000";
end if;
if pc = 4216 then
	inst <= x"44242000";
end if;
if pc = 4220 then
	inst <= x"820010D0";
end if;
if pc = 4224 then
	inst <= x"44262000";
end if;
if pc = 4228 then
	inst <= x"C84000A8";
end if;
if pc = 4232 then
	inst <= x"C86000A4";
end if;
if pc = 4236 then
	inst <= x"48662000";
end if;
if pc = 4240 then
	inst <= x"48662000";
end if;
if pc = 4244 then
	inst <= x"44446000";
end if;
if pc = 4248 then
	inst <= x"C86000A0";
end if;
if pc = 4252 then
	inst <= x"48662000";
end if;
if pc = 4256 then
	inst <= x"48662000";
end if;
if pc = 4260 then
	inst <= x"48662000";
end if;
if pc = 4264 then
	inst <= x"48662000";
end if;
if pc = 4268 then
	inst <= x"40446000";
end if;
if pc = 4272 then
	inst <= x"C860009C";
end if;
if pc = 4276 then
	inst <= x"48662000";
end if;
if pc = 4280 then
	inst <= x"48662000";
end if;
if pc = 4284 then
	inst <= x"48662000";
end if;
if pc = 4288 then
	inst <= x"48662000";
end if;
if pc = 4292 then
	inst <= x"48662000";
end if;
if pc = 4296 then
	inst <= x"48262000";
end if;
if pc = 4300 then
	inst <= x"44242000";
end if;
if pc = 4304 then
	inst <= x"44202000";
end if;
if pc = 4308 then
	inst <= x"C1FDFFFC";
end if;
if pc = 4312 then
	inst <= x"C84000C0";
end if;
if pc = 4316 then
	inst <= x"C86000BC";
end if;
if pc = 4320 then
	inst <= x"C88000B8";
end if;
if pc = 4324 then
	inst <= x"8E24110C";
end if;
if pc = 4328 then
	inst <= x"44224000";
end if;
if pc = 4332 then
	inst <= x"02200001";
end if;
if pc = 4336 then
	inst <= x"C17DFFFC";
end if;
if pc = 4340 then
	inst <= x"03DC0008";
end if;
if pc = 4344 then
	inst <= x"037E000C";
end if;
if pc = 4348 then
	inst <= x"C57DFFFC";
end if;
if pc = 4352 then
	inst <= x"8200084C";
end if;
if pc = 4356 then
	inst <= x"07DC0008";
end if;
if pc = 4360 then
	inst <= x"8200126C";
end if;
if pc = 4364 then
	inst <= x"8E2611C0";
end if;
if pc = 4368 then
	inst <= x"8E82116C";
end if;
if pc = 4372 then
	inst <= x"C84000B4";
end if;
if pc = 4376 then
	inst <= x"48442000";
end if;
if pc = 4380 then
	inst <= x"48442000";
end if;
if pc = 4384 then
	inst <= x"48442000";
end if;
if pc = 4388 then
	inst <= x"44424000";
end if;
if pc = 4392 then
	inst <= x"C86000B0";
end if;
if pc = 4396 then
	inst <= x"48662000";
end if;
if pc = 4400 then
	inst <= x"48662000";
end if;
if pc = 4404 then
	inst <= x"48662000";
end if;
if pc = 4408 then
	inst <= x"48662000";
end if;
if pc = 4412 then
	inst <= x"48662000";
end if;
if pc = 4416 then
	inst <= x"40446000";
end if;
if pc = 4420 then
	inst <= x"C86000AC";
end if;
if pc = 4424 then
	inst <= x"48662000";
end if;
if pc = 4428 then
	inst <= x"48662000";
end if;
if pc = 4432 then
	inst <= x"48662000";
end if;
if pc = 4436 then
	inst <= x"48662000";
end if;
if pc = 4440 then
	inst <= x"48662000";
end if;
if pc = 4444 then
	inst <= x"48662000";
end if;
if pc = 4448 then
	inst <= x"48262000";
end if;
if pc = 4452 then
	inst <= x"44242000";
end if;
if pc = 4456 then
	inst <= x"820011BC";
end if;
if pc = 4460 then
	inst <= x"44262000";
end if;
if pc = 4464 then
	inst <= x"C84000A8";
end if;
if pc = 4468 then
	inst <= x"C86000A4";
end if;
if pc = 4472 then
	inst <= x"48662000";
end if;
if pc = 4476 then
	inst <= x"48662000";
end if;
if pc = 4480 then
	inst <= x"44446000";
end if;
if pc = 4484 then
	inst <= x"C86000A0";
end if;
if pc = 4488 then
	inst <= x"48662000";
end if;
if pc = 4492 then
	inst <= x"48662000";
end if;
if pc = 4496 then
	inst <= x"48662000";
end if;
if pc = 4500 then
	inst <= x"48662000";
end if;
if pc = 4504 then
	inst <= x"40446000";
end if;
if pc = 4508 then
	inst <= x"C860009C";
end if;
if pc = 4512 then
	inst <= x"48662000";
end if;
if pc = 4516 then
	inst <= x"48662000";
end if;
if pc = 4520 then
	inst <= x"48662000";
end if;
if pc = 4524 then
	inst <= x"48662000";
end if;
if pc = 4528 then
	inst <= x"48662000";
end if;
if pc = 4532 then
	inst <= x"48262000";
end if;
if pc = 4536 then
	inst <= x"44242000";
end if;
if pc = 4540 then
	inst <= x"8200126C";
end if;
if pc = 4544 then
	inst <= x"8E82121C";
end if;
if pc = 4548 then
	inst <= x"C84000B4";
end if;
if pc = 4552 then
	inst <= x"48442000";
end if;
if pc = 4556 then
	inst <= x"48442000";
end if;
if pc = 4560 then
	inst <= x"48442000";
end if;
if pc = 4564 then
	inst <= x"44424000";
end if;
if pc = 4568 then
	inst <= x"C86000B0";
end if;
if pc = 4572 then
	inst <= x"48662000";
end if;
if pc = 4576 then
	inst <= x"48662000";
end if;
if pc = 4580 then
	inst <= x"48662000";
end if;
if pc = 4584 then
	inst <= x"48662000";
end if;
if pc = 4588 then
	inst <= x"48662000";
end if;
if pc = 4592 then
	inst <= x"40446000";
end if;
if pc = 4596 then
	inst <= x"C86000AC";
end if;
if pc = 4600 then
	inst <= x"48662000";
end if;
if pc = 4604 then
	inst <= x"48662000";
end if;
if pc = 4608 then
	inst <= x"48662000";
end if;
if pc = 4612 then
	inst <= x"48662000";
end if;
if pc = 4616 then
	inst <= x"48662000";
end if;
if pc = 4620 then
	inst <= x"48662000";
end if;
if pc = 4624 then
	inst <= x"48262000";
end if;
if pc = 4628 then
	inst <= x"44242000";
end if;
if pc = 4632 then
	inst <= x"8200126C";
end if;
if pc = 4636 then
	inst <= x"44262000";
end if;
if pc = 4640 then
	inst <= x"C84000A8";
end if;
if pc = 4644 then
	inst <= x"C86000A4";
end if;
if pc = 4648 then
	inst <= x"48662000";
end if;
if pc = 4652 then
	inst <= x"48662000";
end if;
if pc = 4656 then
	inst <= x"44446000";
end if;
if pc = 4660 then
	inst <= x"C86000A0";
end if;
if pc = 4664 then
	inst <= x"48662000";
end if;
if pc = 4668 then
	inst <= x"48662000";
end if;
if pc = 4672 then
	inst <= x"48662000";
end if;
if pc = 4676 then
	inst <= x"48662000";
end if;
if pc = 4680 then
	inst <= x"40446000";
end if;
if pc = 4684 then
	inst <= x"C860009C";
end if;
if pc = 4688 then
	inst <= x"48662000";
end if;
if pc = 4692 then
	inst <= x"48662000";
end if;
if pc = 4696 then
	inst <= x"48662000";
end if;
if pc = 4700 then
	inst <= x"48662000";
end if;
if pc = 4704 then
	inst <= x"48662000";
end if;
if pc = 4708 then
	inst <= x"48262000";
end if;
if pc = 4712 then
	inst <= x"44242000";
end if;
if pc = 4716 then
	inst <= x"C1FDFFFC";
end if;
if pc = 4720 then
	inst <= x"C8400098";
end if;
if pc = 4724 then
	inst <= x"8E2412AC";
end if;
if pc = 4728 then
	inst <= x"44224000";
end if;
if pc = 4732 then
	inst <= x"8E241288";
end if;
if pc = 4736 then
	inst <= x"44224000";
end if;
if pc = 4740 then
	inst <= x"82001270";
end if;
if pc = 4744 then
	inst <= x"8E0212A4";
end if;
if pc = 4748 then
	inst <= x"C8600090";
end if;
if pc = 4752 then
	inst <= x"8E62129C";
end if;
if pc = 4756 then
	inst <= x"40224000";
end if;
if pc = 4760 then
	inst <= x"82001270";
end if;
if pc = 4764 then
	inst <= x"02200001";
end if;
if pc = 4768 then
	inst <= x"82000B88";
end if;
if pc = 4772 then
	inst <= x"0220FFFF";
end if;
if pc = 4776 then
	inst <= x"82000B88";
end if;
if pc = 4780 then
	inst <= x"8E021484";
end if;
if pc = 4784 then
	inst <= x"C8600090";
end if;
if pc = 4788 then
	inst <= x"8E6212E8";
end if;
if pc = 4792 then
	inst <= x"40224000";
end if;
if pc = 4796 then
	inst <= x"8E2412C8";
end if;
if pc = 4800 then
	inst <= x"44224000";
end if;
if pc = 4804 then
	inst <= x"82001270";
end if;
if pc = 4808 then
	inst <= x"8E0212E0";
end if;
if pc = 4812 then
	inst <= x"8E6212D8";
end if;
if pc = 4816 then
	inst <= x"40224000";
end if;
if pc = 4820 then
	inst <= x"82001270";
end if;
if pc = 4824 then
	inst <= x"02200001";
end if;
if pc = 4828 then
	inst <= x"82000B88";
end if;
if pc = 4832 then
	inst <= x"0220FFFF";
end if;
if pc = 4836 then
	inst <= x"82000B88";
end if;
if pc = 4840 then
	inst <= x"C84000C0";
end if;
if pc = 4844 then
	inst <= x"C86000BC";
end if;
if pc = 4848 then
	inst <= x"C88000B8";
end if;
if pc = 4852 then
	inst <= x"8E24131C";
end if;
if pc = 4856 then
	inst <= x"44224000";
end if;
if pc = 4860 then
	inst <= x"0220FFFF";
end if;
if pc = 4864 then
	inst <= x"C17DFFFC";
end if;
if pc = 4868 then
	inst <= x"03DC0008";
end if;
if pc = 4872 then
	inst <= x"037E000C";
end if;
if pc = 4876 then
	inst <= x"C57DFFFC";
end if;
if pc = 4880 then
	inst <= x"8200084C";
end if;
if pc = 4884 then
	inst <= x"07DC0008";
end if;
if pc = 4888 then
	inst <= x"8200147C";
end if;
if pc = 4892 then
	inst <= x"8E2613D0";
end if;
if pc = 4896 then
	inst <= x"8E821374";
end if;
if pc = 4900 then
	inst <= x"C84000A8";
end if;
if pc = 4904 then
	inst <= x"C86000A4";
end if;
if pc = 4908 then
	inst <= x"48662000";
end if;
if pc = 4912 then
	inst <= x"48662000";
end if;
if pc = 4916 then
	inst <= x"44446000";
end if;
if pc = 4920 then
	inst <= x"C86000A0";
end if;
if pc = 4924 then
	inst <= x"48662000";
end if;
if pc = 4928 then
	inst <= x"48662000";
end if;
if pc = 4932 then
	inst <= x"48662000";
end if;
if pc = 4936 then
	inst <= x"48662000";
end if;
if pc = 4940 then
	inst <= x"40446000";
end if;
if pc = 4944 then
	inst <= x"C860009C";
end if;
if pc = 4948 then
	inst <= x"48662000";
end if;
if pc = 4952 then
	inst <= x"48662000";
end if;
if pc = 4956 then
	inst <= x"48662000";
end if;
if pc = 4960 then
	inst <= x"48662000";
end if;
if pc = 4964 then
	inst <= x"48662000";
end if;
if pc = 4968 then
	inst <= x"48262000";
end if;
if pc = 4972 then
	inst <= x"44242000";
end if;
if pc = 4976 then
	inst <= x"820013CC";
end if;
if pc = 4980 then
	inst <= x"44262000";
end if;
if pc = 4984 then
	inst <= x"C84000B4";
end if;
if pc = 4988 then
	inst <= x"48442000";
end if;
if pc = 4992 then
	inst <= x"48442000";
end if;
if pc = 4996 then
	inst <= x"48442000";
end if;
if pc = 5000 then
	inst <= x"44424000";
end if;
if pc = 5004 then
	inst <= x"C86000B0";
end if;
if pc = 5008 then
	inst <= x"48662000";
end if;
if pc = 5012 then
	inst <= x"48662000";
end if;
if pc = 5016 then
	inst <= x"48662000";
end if;
if pc = 5020 then
	inst <= x"48662000";
end if;
if pc = 5024 then
	inst <= x"48662000";
end if;
if pc = 5028 then
	inst <= x"40446000";
end if;
if pc = 5032 then
	inst <= x"C86000AC";
end if;
if pc = 5036 then
	inst <= x"48662000";
end if;
if pc = 5040 then
	inst <= x"48662000";
end if;
if pc = 5044 then
	inst <= x"48662000";
end if;
if pc = 5048 then
	inst <= x"48662000";
end if;
if pc = 5052 then
	inst <= x"48662000";
end if;
if pc = 5056 then
	inst <= x"48662000";
end if;
if pc = 5060 then
	inst <= x"48262000";
end if;
if pc = 5064 then
	inst <= x"44242000";
end if;
if pc = 5068 then
	inst <= x"8200147C";
end if;
if pc = 5072 then
	inst <= x"8E821424";
end if;
if pc = 5076 then
	inst <= x"C84000A8";
end if;
if pc = 5080 then
	inst <= x"C86000A4";
end if;
if pc = 5084 then
	inst <= x"48662000";
end if;
if pc = 5088 then
	inst <= x"48662000";
end if;
if pc = 5092 then
	inst <= x"44446000";
end if;
if pc = 5096 then
	inst <= x"C86000A0";
end if;
if pc = 5100 then
	inst <= x"48662000";
end if;
if pc = 5104 then
	inst <= x"48662000";
end if;
if pc = 5108 then
	inst <= x"48662000";
end if;
if pc = 5112 then
	inst <= x"48662000";
end if;
if pc = 5116 then
	inst <= x"40446000";
end if;
if pc = 5120 then
	inst <= x"C860009C";
end if;
if pc = 5124 then
	inst <= x"48662000";
end if;
if pc = 5128 then
	inst <= x"48662000";
end if;
if pc = 5132 then
	inst <= x"48662000";
end if;
if pc = 5136 then
	inst <= x"48662000";
end if;
if pc = 5140 then
	inst <= x"48662000";
end if;
if pc = 5144 then
	inst <= x"48262000";
end if;
if pc = 5148 then
	inst <= x"44242000";
end if;
if pc = 5152 then
	inst <= x"8200147C";
end if;
if pc = 5156 then
	inst <= x"44262000";
end if;
if pc = 5160 then
	inst <= x"C84000B4";
end if;
if pc = 5164 then
	inst <= x"48442000";
end if;
if pc = 5168 then
	inst <= x"48442000";
end if;
if pc = 5172 then
	inst <= x"48442000";
end if;
if pc = 5176 then
	inst <= x"44424000";
end if;
if pc = 5180 then
	inst <= x"C86000B0";
end if;
if pc = 5184 then
	inst <= x"48662000";
end if;
if pc = 5188 then
	inst <= x"48662000";
end if;
if pc = 5192 then
	inst <= x"48662000";
end if;
if pc = 5196 then
	inst <= x"48662000";
end if;
if pc = 5200 then
	inst <= x"48662000";
end if;
if pc = 5204 then
	inst <= x"40446000";
end if;
if pc = 5208 then
	inst <= x"C86000AC";
end if;
if pc = 5212 then
	inst <= x"48662000";
end if;
if pc = 5216 then
	inst <= x"48662000";
end if;
if pc = 5220 then
	inst <= x"48662000";
end if;
if pc = 5224 then
	inst <= x"48662000";
end if;
if pc = 5228 then
	inst <= x"48662000";
end if;
if pc = 5232 then
	inst <= x"48662000";
end if;
if pc = 5236 then
	inst <= x"48262000";
end if;
if pc = 5240 then
	inst <= x"44242000";
end if;
if pc = 5244 then
	inst <= x"44202000";
end if;
if pc = 5248 then
	inst <= x"C1FDFFFC";
end if;
if pc = 5252 then
	inst <= x"C84000C0";
end if;
if pc = 5256 then
	inst <= x"C86000BC";
end if;
if pc = 5260 then
	inst <= x"C88000B8";
end if;
if pc = 5264 then
	inst <= x"8E2414B8";
end if;
if pc = 5268 then
	inst <= x"44224000";
end if;
if pc = 5272 then
	inst <= x"02200001";
end if;
if pc = 5276 then
	inst <= x"C17DFFFC";
end if;
if pc = 5280 then
	inst <= x"03DC0008";
end if;
if pc = 5284 then
	inst <= x"037E000C";
end if;
if pc = 5288 then
	inst <= x"C57DFFFC";
end if;
if pc = 5292 then
	inst <= x"8200084C";
end if;
if pc = 5296 then
	inst <= x"07DC0008";
end if;
if pc = 5300 then
	inst <= x"82001618";
end if;
if pc = 5304 then
	inst <= x"8E26156C";
end if;
if pc = 5308 then
	inst <= x"8E821510";
end if;
if pc = 5312 then
	inst <= x"C84000A8";
end if;
if pc = 5316 then
	inst <= x"C86000A4";
end if;
if pc = 5320 then
	inst <= x"48662000";
end if;
if pc = 5324 then
	inst <= x"48662000";
end if;
if pc = 5328 then
	inst <= x"44446000";
end if;
if pc = 5332 then
	inst <= x"C86000A0";
end if;
if pc = 5336 then
	inst <= x"48662000";
end if;
if pc = 5340 then
	inst <= x"48662000";
end if;
if pc = 5344 then
	inst <= x"48662000";
end if;
if pc = 5348 then
	inst <= x"48662000";
end if;
if pc = 5352 then
	inst <= x"40446000";
end if;
if pc = 5356 then
	inst <= x"C860009C";
end if;
if pc = 5360 then
	inst <= x"48662000";
end if;
if pc = 5364 then
	inst <= x"48662000";
end if;
if pc = 5368 then
	inst <= x"48662000";
end if;
if pc = 5372 then
	inst <= x"48662000";
end if;
if pc = 5376 then
	inst <= x"48662000";
end if;
if pc = 5380 then
	inst <= x"48262000";
end if;
if pc = 5384 then
	inst <= x"44242000";
end if;
if pc = 5388 then
	inst <= x"82001568";
end if;
if pc = 5392 then
	inst <= x"44262000";
end if;
if pc = 5396 then
	inst <= x"C84000B4";
end if;
if pc = 5400 then
	inst <= x"48442000";
end if;
if pc = 5404 then
	inst <= x"48442000";
end if;
if pc = 5408 then
	inst <= x"48442000";
end if;
if pc = 5412 then
	inst <= x"44424000";
end if;
if pc = 5416 then
	inst <= x"C86000B0";
end if;
if pc = 5420 then
	inst <= x"48662000";
end if;
if pc = 5424 then
	inst <= x"48662000";
end if;
if pc = 5428 then
	inst <= x"48662000";
end if;
if pc = 5432 then
	inst <= x"48662000";
end if;
if pc = 5436 then
	inst <= x"48662000";
end if;
if pc = 5440 then
	inst <= x"40446000";
end if;
if pc = 5444 then
	inst <= x"C86000AC";
end if;
if pc = 5448 then
	inst <= x"48662000";
end if;
if pc = 5452 then
	inst <= x"48662000";
end if;
if pc = 5456 then
	inst <= x"48662000";
end if;
if pc = 5460 then
	inst <= x"48662000";
end if;
if pc = 5464 then
	inst <= x"48662000";
end if;
if pc = 5468 then
	inst <= x"48662000";
end if;
if pc = 5472 then
	inst <= x"48262000";
end if;
if pc = 5476 then
	inst <= x"44242000";
end if;
if pc = 5480 then
	inst <= x"82001618";
end if;
if pc = 5484 then
	inst <= x"8E8215C0";
end if;
if pc = 5488 then
	inst <= x"C84000A8";
end if;
if pc = 5492 then
	inst <= x"C86000A4";
end if;
if pc = 5496 then
	inst <= x"48662000";
end if;
if pc = 5500 then
	inst <= x"48662000";
end if;
if pc = 5504 then
	inst <= x"44446000";
end if;
if pc = 5508 then
	inst <= x"C86000A0";
end if;
if pc = 5512 then
	inst <= x"48662000";
end if;
if pc = 5516 then
	inst <= x"48662000";
end if;
if pc = 5520 then
	inst <= x"48662000";
end if;
if pc = 5524 then
	inst <= x"48662000";
end if;
if pc = 5528 then
	inst <= x"40446000";
end if;
if pc = 5532 then
	inst <= x"C860009C";
end if;
if pc = 5536 then
	inst <= x"48662000";
end if;
if pc = 5540 then
	inst <= x"48662000";
end if;
if pc = 5544 then
	inst <= x"48662000";
end if;
if pc = 5548 then
	inst <= x"48662000";
end if;
if pc = 5552 then
	inst <= x"48662000";
end if;
if pc = 5556 then
	inst <= x"48262000";
end if;
if pc = 5560 then
	inst <= x"44242000";
end if;
if pc = 5564 then
	inst <= x"82001618";
end if;
if pc = 5568 then
	inst <= x"44262000";
end if;
if pc = 5572 then
	inst <= x"C84000B4";
end if;
if pc = 5576 then
	inst <= x"48442000";
end if;
if pc = 5580 then
	inst <= x"48442000";
end if;
if pc = 5584 then
	inst <= x"48442000";
end if;
if pc = 5588 then
	inst <= x"44424000";
end if;
if pc = 5592 then
	inst <= x"C86000B0";
end if;
if pc = 5596 then
	inst <= x"48662000";
end if;
if pc = 5600 then
	inst <= x"48662000";
end if;
if pc = 5604 then
	inst <= x"48662000";
end if;
if pc = 5608 then
	inst <= x"48662000";
end if;
if pc = 5612 then
	inst <= x"48662000";
end if;
if pc = 5616 then
	inst <= x"40446000";
end if;
if pc = 5620 then
	inst <= x"C86000AC";
end if;
if pc = 5624 then
	inst <= x"48662000";
end if;
if pc = 5628 then
	inst <= x"48662000";
end if;
if pc = 5632 then
	inst <= x"48662000";
end if;
if pc = 5636 then
	inst <= x"48662000";
end if;
if pc = 5640 then
	inst <= x"48662000";
end if;
if pc = 5644 then
	inst <= x"48662000";
end if;
if pc = 5648 then
	inst <= x"48262000";
end if;
if pc = 5652 then
	inst <= x"44242000";
end if;
if pc = 5656 then
	inst <= x"C1FDFFFC";
end if;
if pc = 5660 then
	inst <= x"C8220000";
end if;
if pc = 5664 then
	inst <= x"48222000";
end if;
if pc = 5668 then
	inst <= x"C8420004";
end if;
if pc = 5672 then
	inst <= x"48444000";
end if;
if pc = 5676 then
	inst <= x"40224000";
end if;
if pc = 5680 then
	inst <= x"C8420008";
end if;
if pc = 5684 then
	inst <= x"48444000";
end if;
if pc = 5688 then
	inst <= x"40224000";
end if;
if pc = 5692 then
	inst <= x"C43C0000";
end if;
if pc = 5696 then
	inst <= x"C45C0004";
end if;
if pc = 5700 then
	inst <= x"C17DFFFC";
end if;
if pc = 5704 then
	inst <= x"03DC0010";
end if;
if pc = 5708 then
	inst <= x"037E000C";
end if;
if pc = 5712 then
	inst <= x"C57DFFFC";
end if;
if pc = 5716 then
	inst <= x"8200083C";
end if;
if pc = 5720 then
	inst <= x"07DC0010";
end if;
if pc = 5724 then
	inst <= x"8A2016A4";
end if;
if pc = 5728 then
	inst <= x"C03C0004";
end if;
if pc = 5732 then
	inst <= x"82201688";
end if;
if pc = 5736 then
	inst <= x"C17DFFFC";
end if;
if pc = 5740 then
	inst <= x"03DC0010";
end if;
if pc = 5744 then
	inst <= x"037E000C";
end if;
if pc = 5748 then
	inst <= x"C57DFFFC";
end if;
if pc = 5752 then
	inst <= x"82000844";
end if;
if pc = 5756 then
	inst <= x"07DC0010";
end if;
if pc = 5760 then
	inst <= x"44202000";
end if;
if pc = 5764 then
	inst <= x"820016A0";
end if;
if pc = 5768 then
	inst <= x"C17DFFFC";
end if;
if pc = 5772 then
	inst <= x"03DC0010";
end if;
if pc = 5776 then
	inst <= x"037E000C";
end if;
if pc = 5780 then
	inst <= x"C57DFFFC";
end if;
if pc = 5784 then
	inst <= x"82000844";
end if;
if pc = 5788 then
	inst <= x"07DC0010";
end if;
if pc = 5792 then
	inst <= x"820016A8";
end if;
if pc = 5796 then
	inst <= x"C82000A8";
end if;
if pc = 5800 then
	inst <= x"C03C0000";
end if;
if pc = 5804 then
	inst <= x"C8420000";
end if;
if pc = 5808 then
	inst <= x"48442000";
end if;
if pc = 5812 then
	inst <= x"CC420000";
end if;
if pc = 5816 then
	inst <= x"C8420004";
end if;
if pc = 5820 then
	inst <= x"48442000";
end if;
if pc = 5824 then
	inst <= x"CC420004";
end if;
if pc = 5828 then
	inst <= x"C8420008";
end if;
if pc = 5832 then
	inst <= x"48242000";
end if;
if pc = 5836 then
	inst <= x"CC220008";
end if;
if pc = 5840 then
	inst <= x"C1FDFFFC";
end if;
if pc = 5844 then
	inst <= x"022001B8";
end if;
if pc = 5848 then
	inst <= x"C43C0000";
end if;
if pc = 5852 then
	inst <= x"C17DFFFC";
end if;
if pc = 5856 then
	inst <= x"03DC000C";
end if;
if pc = 5860 then
	inst <= x"037E000C";
end if;
if pc = 5864 then
	inst <= x"C57DFFFC";
end if;
if pc = 5868 then
	inst <= x"820007C0";
end if;
if pc = 5872 then
	inst <= x"07DC000C";
end if;
if pc = 5876 then
	inst <= x"C03C0000";
end if;
if pc = 5880 then
	inst <= x"CC220000";
end if;
if pc = 5884 then
	inst <= x"C17DFFFC";
end if;
if pc = 5888 then
	inst <= x"03DC000C";
end if;
if pc = 5892 then
	inst <= x"037E000C";
end if;
if pc = 5896 then
	inst <= x"C57DFFFC";
end if;
if pc = 5900 then
	inst <= x"820007C0";
end if;
if pc = 5904 then
	inst <= x"07DC000C";
end if;
if pc = 5908 then
	inst <= x"C03C0000";
end if;
if pc = 5912 then
	inst <= x"CC220004";
end if;
if pc = 5916 then
	inst <= x"C17DFFFC";
end if;
if pc = 5920 then
	inst <= x"03DC000C";
end if;
if pc = 5924 then
	inst <= x"037E000C";
end if;
if pc = 5928 then
	inst <= x"C57DFFFC";
end if;
if pc = 5932 then
	inst <= x"820007C0";
end if;
if pc = 5936 then
	inst <= x"07DC000C";
end if;
if pc = 5940 then
	inst <= x"C03C0000";
end if;
if pc = 5944 then
	inst <= x"CC220008";
end if;
if pc = 5948 then
	inst <= x"C17DFFFC";
end if;
if pc = 5952 then
	inst <= x"03DC000C";
end if;
if pc = 5956 then
	inst <= x"037E000C";
end if;
if pc = 5960 then
	inst <= x"C57DFFFC";
end if;
if pc = 5964 then
	inst <= x"820007C0";
end if;
if pc = 5968 then
	inst <= x"07DC000C";
end if;
if pc = 5972 then
	inst <= x"C840008C";
end if;
if pc = 5976 then
	inst <= x"48224000";
end if;
if pc = 5980 then
	inst <= x"C8600098";
end if;
if pc = 5984 then
	inst <= x"CC5C0008";
end if;
if pc = 5988 then
	inst <= x"CC7C0010";
end if;
if pc = 5992 then
	inst <= x"CC3C0018";
end if;
if pc = 5996 then
	inst <= x"8E261794";
end if;
if pc = 6000 then
	inst <= x"44826000";
end if;
if pc = 6004 then
	inst <= x"C17DFFFC";
end if;
if pc = 6008 then
	inst <= x"40208000";
end if;
if pc = 6012 then
	inst <= x"03DC0028";
end if;
if pc = 6016 then
	inst <= x"037E000C";
end if;
if pc = 6020 then
	inst <= x"C57DFFFC";
end if;
if pc = 6024 then
	inst <= x"82001270";
end if;
if pc = 6028 then
	inst <= x"07DC0028";
end if;
if pc = 6032 then
	inst <= x"82001800";
end if;
if pc = 6036 then
	inst <= x"8E0217E4";
end if;
if pc = 6040 then
	inst <= x"C8800090";
end if;
if pc = 6044 then
	inst <= x"8E8217C4";
end if;
if pc = 6048 then
	inst <= x"40826000";
end if;
if pc = 6052 then
	inst <= x"C17DFFFC";
end if;
if pc = 6056 then
	inst <= x"40208000";
end if;
if pc = 6060 then
	inst <= x"03DC0028";
end if;
if pc = 6064 then
	inst <= x"037E000C";
end if;
if pc = 6068 then
	inst <= x"C57DFFFC";
end if;
if pc = 6072 then
	inst <= x"82001270";
end if;
if pc = 6076 then
	inst <= x"07DC0028";
end if;
if pc = 6080 then
	inst <= x"820017E0";
end if;
if pc = 6084 then
	inst <= x"02200001";
end if;
if pc = 6088 then
	inst <= x"C17DFFFC";
end if;
if pc = 6092 then
	inst <= x"03DC0028";
end if;
if pc = 6096 then
	inst <= x"037E000C";
end if;
if pc = 6100 then
	inst <= x"C57DFFFC";
end if;
if pc = 6104 then
	inst <= x"82000B88";
end if;
if pc = 6108 then
	inst <= x"07DC0028";
end if;
if pc = 6112 then
	inst <= x"82001800";
end if;
if pc = 6116 then
	inst <= x"0220FFFF";
end if;
if pc = 6120 then
	inst <= x"C17DFFFC";
end if;
if pc = 6124 then
	inst <= x"03DC0028";
end if;
if pc = 6128 then
	inst <= x"037E000C";
end if;
if pc = 6132 then
	inst <= x"C57DFFFC";
end if;
if pc = 6136 then
	inst <= x"82000B88";
end if;
if pc = 6140 then
	inst <= x"07DC0028";
end if;
if pc = 6144 then
	inst <= x"C85C0010";
end if;
if pc = 6148 then
	inst <= x"C87C0018";
end if;
if pc = 6152 then
	inst <= x"CC3C0020";
end if;
if pc = 6156 then
	inst <= x"8E641834";
end if;
if pc = 6160 then
	inst <= x"44664000";
end if;
if pc = 6164 then
	inst <= x"C17DFFFC";
end if;
if pc = 6168 then
	inst <= x"40206000";
end if;
if pc = 6172 then
	inst <= x"03DC0030";
end if;
if pc = 6176 then
	inst <= x"037E000C";
end if;
if pc = 6180 then
	inst <= x"C57DFFFC";
end if;
if pc = 6184 then
	inst <= x"82000EC4";
end if;
if pc = 6188 then
	inst <= x"07DC0030";
end if;
if pc = 6192 then
	inst <= x"820018A8";
end if;
if pc = 6196 then
	inst <= x"8E061888";
end if;
if pc = 6200 then
	inst <= x"C8800090";
end if;
if pc = 6204 then
	inst <= x"8E861864";
end if;
if pc = 6208 then
	inst <= x"40664000";
end if;
if pc = 6212 then
	inst <= x"C17DFFFC";
end if;
if pc = 6216 then
	inst <= x"40206000";
end if;
if pc = 6220 then
	inst <= x"03DC0030";
end if;
if pc = 6224 then
	inst <= x"037E000C";
end if;
if pc = 6228 then
	inst <= x"C57DFFFC";
end if;
if pc = 6232 then
	inst <= x"82000EC4";
end if;
if pc = 6236 then
	inst <= x"07DC0030";
end if;
if pc = 6240 then
	inst <= x"82001884";
end if;
if pc = 6244 then
	inst <= x"02200001";
end if;
if pc = 6248 then
	inst <= x"C17DFFFC";
end if;
if pc = 6252 then
	inst <= x"40206000";
end if;
if pc = 6256 then
	inst <= x"03DC0030";
end if;
if pc = 6260 then
	inst <= x"037E000C";
end if;
if pc = 6264 then
	inst <= x"C57DFFFC";
end if;
if pc = 6268 then
	inst <= x"8200084C";
end if;
if pc = 6272 then
	inst <= x"07DC0030";
end if;
if pc = 6276 then
	inst <= x"820018A8";
end if;
if pc = 6280 then
	inst <= x"0220FFFF";
end if;
if pc = 6284 then
	inst <= x"C17DFFFC";
end if;
if pc = 6288 then
	inst <= x"40206000";
end if;
if pc = 6292 then
	inst <= x"03DC0030";
end if;
if pc = 6296 then
	inst <= x"037E000C";
end if;
if pc = 6300 then
	inst <= x"C57DFFFC";
end if;
if pc = 6304 then
	inst <= x"8200084C";
end if;
if pc = 6308 then
	inst <= x"07DC0030";
end if;
if pc = 6312 then
	inst <= x"CC3C0028";
end if;
if pc = 6316 then
	inst <= x"C17DFFFC";
end if;
if pc = 6320 then
	inst <= x"03DC0038";
end if;
if pc = 6324 then
	inst <= x"037E000C";
end if;
if pc = 6328 then
	inst <= x"C57DFFFC";
end if;
if pc = 6332 then
	inst <= x"820007C0";
end if;
if pc = 6336 then
	inst <= x"07DC0038";
end if;
if pc = 6340 then
	inst <= x"C85C0008";
end if;
if pc = 6344 then
	inst <= x"48224000";
end if;
if pc = 6348 then
	inst <= x"C85C0010";
end if;
if pc = 6352 then
	inst <= x"CC3C0030";
end if;
if pc = 6356 then
	inst <= x"8E2418FC";
end if;
if pc = 6360 then
	inst <= x"44624000";
end if;
if pc = 6364 then
	inst <= x"C17DFFFC";
end if;
if pc = 6368 then
	inst <= x"40206000";
end if;
if pc = 6372 then
	inst <= x"03DC0040";
end if;
if pc = 6376 then
	inst <= x"037E000C";
end if;
if pc = 6380 then
	inst <= x"C57DFFFC";
end if;
if pc = 6384 then
	inst <= x"82001270";
end if;
if pc = 6388 then
	inst <= x"07DC0040";
end if;
if pc = 6392 then
	inst <= x"82001968";
end if;
if pc = 6396 then
	inst <= x"8E02194C";
end if;
if pc = 6400 then
	inst <= x"C8600090";
end if;
if pc = 6404 then
	inst <= x"8E62192C";
end if;
if pc = 6408 then
	inst <= x"40624000";
end if;
if pc = 6412 then
	inst <= x"C17DFFFC";
end if;
if pc = 6416 then
	inst <= x"40206000";
end if;
if pc = 6420 then
	inst <= x"03DC0040";
end if;
if pc = 6424 then
	inst <= x"037E000C";
end if;
if pc = 6428 then
	inst <= x"C57DFFFC";
end if;
if pc = 6432 then
	inst <= x"82001270";
end if;
if pc = 6436 then
	inst <= x"07DC0040";
end if;
if pc = 6440 then
	inst <= x"82001948";
end if;
if pc = 6444 then
	inst <= x"02200001";
end if;
if pc = 6448 then
	inst <= x"C17DFFFC";
end if;
if pc = 6452 then
	inst <= x"03DC0040";
end if;
if pc = 6456 then
	inst <= x"037E000C";
end if;
if pc = 6460 then
	inst <= x"C57DFFFC";
end if;
if pc = 6464 then
	inst <= x"82000B88";
end if;
if pc = 6468 then
	inst <= x"07DC0040";
end if;
if pc = 6472 then
	inst <= x"82001968";
end if;
if pc = 6476 then
	inst <= x"0220FFFF";
end if;
if pc = 6480 then
	inst <= x"C17DFFFC";
end if;
if pc = 6484 then
	inst <= x"03DC0040";
end if;
if pc = 6488 then
	inst <= x"037E000C";
end if;
if pc = 6492 then
	inst <= x"C57DFFFC";
end if;
if pc = 6496 then
	inst <= x"82000B88";
end if;
if pc = 6500 then
	inst <= x"07DC0040";
end if;
if pc = 6504 then
	inst <= x"C85C0010";
end if;
if pc = 6508 then
	inst <= x"C87C0030";
end if;
if pc = 6512 then
	inst <= x"CC3C0038";
end if;
if pc = 6516 then
	inst <= x"8E64199C";
end if;
if pc = 6520 then
	inst <= x"44464000";
end if;
if pc = 6524 then
	inst <= x"C17DFFFC";
end if;
if pc = 6528 then
	inst <= x"40204000";
end if;
if pc = 6532 then
	inst <= x"03DC0048";
end if;
if pc = 6536 then
	inst <= x"037E000C";
end if;
if pc = 6540 then
	inst <= x"C57DFFFC";
end if;
if pc = 6544 then
	inst <= x"82000EC4";
end if;
if pc = 6548 then
	inst <= x"07DC0048";
end if;
if pc = 6552 then
	inst <= x"82001A10";
end if;
if pc = 6556 then
	inst <= x"8E0619F0";
end if;
if pc = 6560 then
	inst <= x"C8800090";
end if;
if pc = 6564 then
	inst <= x"8E8619CC";
end if;
if pc = 6568 then
	inst <= x"40464000";
end if;
if pc = 6572 then
	inst <= x"C17DFFFC";
end if;
if pc = 6576 then
	inst <= x"40204000";
end if;
if pc = 6580 then
	inst <= x"03DC0048";
end if;
if pc = 6584 then
	inst <= x"037E000C";
end if;
if pc = 6588 then
	inst <= x"C57DFFFC";
end if;
if pc = 6592 then
	inst <= x"82000EC4";
end if;
if pc = 6596 then
	inst <= x"07DC0048";
end if;
if pc = 6600 then
	inst <= x"820019EC";
end if;
if pc = 6604 then
	inst <= x"02200001";
end if;
if pc = 6608 then
	inst <= x"C17DFFFC";
end if;
if pc = 6612 then
	inst <= x"40206000";
end if;
if pc = 6616 then
	inst <= x"03DC0048";
end if;
if pc = 6620 then
	inst <= x"037E000C";
end if;
if pc = 6624 then
	inst <= x"C57DFFFC";
end if;
if pc = 6628 then
	inst <= x"8200084C";
end if;
if pc = 6632 then
	inst <= x"07DC0048";
end if;
if pc = 6636 then
	inst <= x"82001A10";
end if;
if pc = 6640 then
	inst <= x"0220FFFF";
end if;
if pc = 6644 then
	inst <= x"C17DFFFC";
end if;
if pc = 6648 then
	inst <= x"40206000";
end if;
if pc = 6652 then
	inst <= x"03DC0048";
end if;
if pc = 6656 then
	inst <= x"037E000C";
end if;
if pc = 6660 then
	inst <= x"C57DFFFC";
end if;
if pc = 6664 then
	inst <= x"8200084C";
end if;
if pc = 6668 then
	inst <= x"07DC0048";
end if;
if pc = 6672 then
	inst <= x"0220033C";
end if;
if pc = 6676 then
	inst <= x"C85C0020";
end if;
if pc = 6680 then
	inst <= x"48642000";
end if;
if pc = 6684 then
	inst <= x"C8800088";
end if;
if pc = 6688 then
	inst <= x"48668000";
end if;
if pc = 6692 then
	inst <= x"CC620000";
end if;
if pc = 6696 then
	inst <= x"C8600084";
end if;
if pc = 6700 then
	inst <= x"C8BC0028";
end if;
if pc = 6704 then
	inst <= x"486A6000";
end if;
if pc = 6708 then
	inst <= x"CC620004";
end if;
if pc = 6712 then
	inst <= x"C87C0038";
end if;
if pc = 6716 then
	inst <= x"48C46000";
end if;
if pc = 6720 then
	inst <= x"488C8000";
end if;
if pc = 6724 then
	inst <= x"CC820008";
end if;
if pc = 6728 then
	inst <= x"02400324";
end if;
if pc = 6732 then
	inst <= x"CC640000";
end if;
if pc = 6736 then
	inst <= x"CC040004";
end if;
if pc = 6740 then
	inst <= x"44802000";
end if;
if pc = 6744 then
	inst <= x"CC840008";
end if;
if pc = 6748 then
	inst <= x"02400330";
end if;
if pc = 6752 then
	inst <= x"4480A000";
end if;
if pc = 6756 then
	inst <= x"48282000";
end if;
if pc = 6760 then
	inst <= x"CC240000";
end if;
if pc = 6764 then
	inst <= x"44204000";
end if;
if pc = 6768 then
	inst <= x"CC240004";
end if;
if pc = 6772 then
	inst <= x"48286000";
end if;
if pc = 6776 then
	inst <= x"CC240008";
end if;
if pc = 6780 then
	inst <= x"024001C4";
end if;
if pc = 6784 then
	inst <= x"C07C0000";
end if;
if pc = 6788 then
	inst <= x"C8260000";
end if;
if pc = 6792 then
	inst <= x"C8420000";
end if;
if pc = 6796 then
	inst <= x"44224000";
end if;
if pc = 6800 then
	inst <= x"CC240000";
end if;
if pc = 6804 then
	inst <= x"C8260004";
end if;
if pc = 6808 then
	inst <= x"C8420004";
end if;
if pc = 6812 then
	inst <= x"44224000";
end if;
if pc = 6816 then
	inst <= x"CC240004";
end if;
if pc = 6820 then
	inst <= x"C8260008";
end if;
if pc = 6824 then
	inst <= x"C8420008";
end if;
if pc = 6828 then
	inst <= x"44224000";
end if;
if pc = 6832 then
	inst <= x"CC240008";
end if;
if pc = 6836 then
	inst <= x"C1FDFFFC";
end if;
if pc = 6840 then
	inst <= x"C17DFFFC";
end if;
if pc = 6844 then
	inst <= x"03DC0008";
end if;
if pc = 6848 then
	inst <= x"037E000C";
end if;
if pc = 6852 then
	inst <= x"C57DFFFC";
end if;
if pc = 6856 then
	inst <= x"82000794";
end if;
if pc = 6860 then
	inst <= x"07DC0008";
end if;
if pc = 6864 then
	inst <= x"C17DFFFC";
end if;
if pc = 6868 then
	inst <= x"03DC0008";
end if;
if pc = 6872 then
	inst <= x"037E000C";
end if;
if pc = 6876 then
	inst <= x"C57DFFFC";
end if;
if pc = 6880 then
	inst <= x"820007C0";
end if;
if pc = 6884 then
	inst <= x"07DC0008";
end if;
if pc = 6888 then
	inst <= x"C840008C";
end if;
if pc = 6892 then
	inst <= x"48224000";
end if;
if pc = 6896 then
	inst <= x"C8600098";
end if;
if pc = 6900 then
	inst <= x"CC7C0000";
end if;
if pc = 6904 then
	inst <= x"CC3C0008";
end if;
if pc = 6908 then
	inst <= x"CC5C0010";
end if;
if pc = 6912 then
	inst <= x"8E261B28";
end if;
if pc = 6916 then
	inst <= x"44826000";
end if;
if pc = 6920 then
	inst <= x"C17DFFFC";
end if;
if pc = 6924 then
	inst <= x"40208000";
end if;
if pc = 6928 then
	inst <= x"03DC0020";
end if;
if pc = 6932 then
	inst <= x"037E000C";
end if;
if pc = 6936 then
	inst <= x"C57DFFFC";
end if;
if pc = 6940 then
	inst <= x"82000EC4";
end if;
if pc = 6944 then
	inst <= x"07DC0020";
end if;
if pc = 6948 then
	inst <= x"82001B94";
end if;
if pc = 6952 then
	inst <= x"8E021B78";
end if;
if pc = 6956 then
	inst <= x"C8800090";
end if;
if pc = 6960 then
	inst <= x"8E821B58";
end if;
if pc = 6964 then
	inst <= x"40826000";
end if;
if pc = 6968 then
	inst <= x"C17DFFFC";
end if;
if pc = 6972 then
	inst <= x"40208000";
end if;
if pc = 6976 then
	inst <= x"03DC0020";
end if;
if pc = 6980 then
	inst <= x"037E000C";
end if;
if pc = 6984 then
	inst <= x"C57DFFFC";
end if;
if pc = 6988 then
	inst <= x"82000EC4";
end if;
if pc = 6992 then
	inst <= x"07DC0020";
end if;
if pc = 6996 then
	inst <= x"82001B74";
end if;
if pc = 7000 then
	inst <= x"02200001";
end if;
if pc = 7004 then
	inst <= x"C17DFFFC";
end if;
if pc = 7008 then
	inst <= x"03DC0020";
end if;
if pc = 7012 then
	inst <= x"037E000C";
end if;
if pc = 7016 then
	inst <= x"C57DFFFC";
end if;
if pc = 7020 then
	inst <= x"8200084C";
end if;
if pc = 7024 then
	inst <= x"07DC0020";
end if;
if pc = 7028 then
	inst <= x"82001B94";
end if;
if pc = 7032 then
	inst <= x"0220FFFF";
end if;
if pc = 7036 then
	inst <= x"C17DFFFC";
end if;
if pc = 7040 then
	inst <= x"03DC0020";
end if;
if pc = 7044 then
	inst <= x"037E000C";
end if;
if pc = 7048 then
	inst <= x"C57DFFFC";
end if;
if pc = 7052 then
	inst <= x"8200084C";
end if;
if pc = 7056 then
	inst <= x"07DC0020";
end if;
if pc = 7060 then
	inst <= x"022001D0";
end if;
if pc = 7064 then
	inst <= x"44202000";
end if;
if pc = 7068 then
	inst <= x"CC220004";
end if;
if pc = 7072 then
	inst <= x"C43C0018";
end if;
if pc = 7076 then
	inst <= x"C17DFFFC";
end if;
if pc = 7080 then
	inst <= x"03DC0024";
end if;
if pc = 7084 then
	inst <= x"037E000C";
end if;
if pc = 7088 then
	inst <= x"C57DFFFC";
end if;
if pc = 7092 then
	inst <= x"820007C0";
end if;
if pc = 7096 then
	inst <= x"07DC0024";
end if;
if pc = 7100 then
	inst <= x"C85C0010";
end if;
if pc = 7104 then
	inst <= x"48224000";
end if;
if pc = 7108 then
	inst <= x"C85C0000";
end if;
if pc = 7112 then
	inst <= x"C87C0008";
end if;
if pc = 7116 then
	inst <= x"CC3C0020";
end if;
if pc = 7120 then
	inst <= x"8E641BF8";
end if;
if pc = 7124 then
	inst <= x"44664000";
end if;
if pc = 7128 then
	inst <= x"C17DFFFC";
end if;
if pc = 7132 then
	inst <= x"40206000";
end if;
if pc = 7136 then
	inst <= x"03DC0030";
end if;
if pc = 7140 then
	inst <= x"037E000C";
end if;
if pc = 7144 then
	inst <= x"C57DFFFC";
end if;
if pc = 7148 then
	inst <= x"82001270";
end if;
if pc = 7152 then
	inst <= x"07DC0030";
end if;
if pc = 7156 then
	inst <= x"82001C6C";
end if;
if pc = 7160 then
	inst <= x"8E061C4C";
end if;
if pc = 7164 then
	inst <= x"C8800090";
end if;
if pc = 7168 then
	inst <= x"8E861C28";
end if;
if pc = 7172 then
	inst <= x"40664000";
end if;
if pc = 7176 then
	inst <= x"C17DFFFC";
end if;
if pc = 7180 then
	inst <= x"40206000";
end if;
if pc = 7184 then
	inst <= x"03DC0030";
end if;
if pc = 7188 then
	inst <= x"037E000C";
end if;
if pc = 7192 then
	inst <= x"C57DFFFC";
end if;
if pc = 7196 then
	inst <= x"82001270";
end if;
if pc = 7200 then
	inst <= x"07DC0030";
end if;
if pc = 7204 then
	inst <= x"82001C48";
end if;
if pc = 7208 then
	inst <= x"02200001";
end if;
if pc = 7212 then
	inst <= x"C17DFFFC";
end if;
if pc = 7216 then
	inst <= x"40206000";
end if;
if pc = 7220 then
	inst <= x"03DC0030";
end if;
if pc = 7224 then
	inst <= x"037E000C";
end if;
if pc = 7228 then
	inst <= x"C57DFFFC";
end if;
if pc = 7232 then
	inst <= x"82000B88";
end if;
if pc = 7236 then
	inst <= x"07DC0030";
end if;
if pc = 7240 then
	inst <= x"82001C6C";
end if;
if pc = 7244 then
	inst <= x"0220FFFF";
end if;
if pc = 7248 then
	inst <= x"C17DFFFC";
end if;
if pc = 7252 then
	inst <= x"40206000";
end if;
if pc = 7256 then
	inst <= x"03DC0030";
end if;
if pc = 7260 then
	inst <= x"037E000C";
end if;
if pc = 7264 then
	inst <= x"C57DFFFC";
end if;
if pc = 7268 then
	inst <= x"82000B88";
end if;
if pc = 7272 then
	inst <= x"07DC0030";
end if;
if pc = 7276 then
	inst <= x"C85C0000";
end if;
if pc = 7280 then
	inst <= x"C87C0020";
end if;
if pc = 7284 then
	inst <= x"CC3C0028";
end if;
if pc = 7288 then
	inst <= x"8E641CA0";
end if;
if pc = 7292 then
	inst <= x"44864000";
end if;
if pc = 7296 then
	inst <= x"C17DFFFC";
end if;
if pc = 7300 then
	inst <= x"40208000";
end if;
if pc = 7304 then
	inst <= x"03DC0038";
end if;
if pc = 7308 then
	inst <= x"037E000C";
end if;
if pc = 7312 then
	inst <= x"C57DFFFC";
end if;
if pc = 7316 then
	inst <= x"82000EC4";
end if;
if pc = 7320 then
	inst <= x"07DC0038";
end if;
if pc = 7324 then
	inst <= x"82001D14";
end if;
if pc = 7328 then
	inst <= x"8E061CF4";
end if;
if pc = 7332 then
	inst <= x"C8800090";
end if;
if pc = 7336 then
	inst <= x"8E861CD0";
end if;
if pc = 7340 then
	inst <= x"40864000";
end if;
if pc = 7344 then
	inst <= x"C17DFFFC";
end if;
if pc = 7348 then
	inst <= x"40208000";
end if;
if pc = 7352 then
	inst <= x"03DC0038";
end if;
if pc = 7356 then
	inst <= x"037E000C";
end if;
if pc = 7360 then
	inst <= x"C57DFFFC";
end if;
if pc = 7364 then
	inst <= x"82000EC4";
end if;
if pc = 7368 then
	inst <= x"07DC0038";
end if;
if pc = 7372 then
	inst <= x"82001CF0";
end if;
if pc = 7376 then
	inst <= x"02200001";
end if;
if pc = 7380 then
	inst <= x"C17DFFFC";
end if;
if pc = 7384 then
	inst <= x"40206000";
end if;
if pc = 7388 then
	inst <= x"03DC0038";
end if;
if pc = 7392 then
	inst <= x"037E000C";
end if;
if pc = 7396 then
	inst <= x"C57DFFFC";
end if;
if pc = 7400 then
	inst <= x"8200084C";
end if;
if pc = 7404 then
	inst <= x"07DC0038";
end if;
if pc = 7408 then
	inst <= x"82001D14";
end if;
if pc = 7412 then
	inst <= x"0220FFFF";
end if;
if pc = 7416 then
	inst <= x"C17DFFFC";
end if;
if pc = 7420 then
	inst <= x"40206000";
end if;
if pc = 7424 then
	inst <= x"03DC0038";
end if;
if pc = 7428 then
	inst <= x"037E000C";
end if;
if pc = 7432 then
	inst <= x"C57DFFFC";
end if;
if pc = 7436 then
	inst <= x"8200084C";
end if;
if pc = 7440 then
	inst <= x"07DC0038";
end if;
if pc = 7444 then
	inst <= x"C85C0028";
end if;
if pc = 7448 then
	inst <= x"48242000";
end if;
if pc = 7452 then
	inst <= x"C03C0018";
end if;
if pc = 7456 then
	inst <= x"CC220000";
end if;
if pc = 7460 then
	inst <= x"C83C0000";
end if;
if pc = 7464 then
	inst <= x"C87C0020";
end if;
if pc = 7468 then
	inst <= x"8E621D50";
end if;
if pc = 7472 then
	inst <= x"44262000";
end if;
if pc = 7476 then
	inst <= x"C17DFFFC";
end if;
if pc = 7480 then
	inst <= x"03DC0038";
end if;
if pc = 7484 then
	inst <= x"037E000C";
end if;
if pc = 7488 then
	inst <= x"C57DFFFC";
end if;
if pc = 7492 then
	inst <= x"82001270";
end if;
if pc = 7496 then
	inst <= x"07DC0038";
end if;
if pc = 7500 then
	inst <= x"82001DC8";
end if;
if pc = 7504 then
	inst <= x"8E061DA4";
end if;
if pc = 7508 then
	inst <= x"C8800090";
end if;
if pc = 7512 then
	inst <= x"8E861D7C";
end if;
if pc = 7516 then
	inst <= x"40262000";
end if;
if pc = 7520 then
	inst <= x"C17DFFFC";
end if;
if pc = 7524 then
	inst <= x"03DC0038";
end if;
if pc = 7528 then
	inst <= x"037E000C";
end if;
if pc = 7532 then
	inst <= x"C57DFFFC";
end if;
if pc = 7536 then
	inst <= x"82001270";
end if;
if pc = 7540 then
	inst <= x"07DC0038";
end if;
if pc = 7544 then
	inst <= x"82001DA0";
end if;
if pc = 7548 then
	inst <= x"02400001";
end if;
if pc = 7552 then
	inst <= x"C17DFFFC";
end if;
if pc = 7556 then
	inst <= x"00240000";
end if;
if pc = 7560 then
	inst <= x"40206000";
end if;
if pc = 7564 then
	inst <= x"03DC0038";
end if;
if pc = 7568 then
	inst <= x"037E000C";
end if;
if pc = 7572 then
	inst <= x"C57DFFFC";
end if;
if pc = 7576 then
	inst <= x"82000B88";
end if;
if pc = 7580 then
	inst <= x"07DC0038";
end if;
if pc = 7584 then
	inst <= x"82001DC8";
end if;
if pc = 7588 then
	inst <= x"0240FFFF";
end if;
if pc = 7592 then
	inst <= x"C17DFFFC";
end if;
if pc = 7596 then
	inst <= x"00240000";
end if;
if pc = 7600 then
	inst <= x"40206000";
end if;
if pc = 7604 then
	inst <= x"03DC0038";
end if;
if pc = 7608 then
	inst <= x"037E000C";
end if;
if pc = 7612 then
	inst <= x"C57DFFFC";
end if;
if pc = 7616 then
	inst <= x"82000B88";
end if;
if pc = 7620 then
	inst <= x"07DC0038";
end if;
if pc = 7624 then
	inst <= x"C85C0028";
end if;
if pc = 7628 then
	inst <= x"48242000";
end if;
if pc = 7632 then
	inst <= x"C03C0018";
end if;
if pc = 7636 then
	inst <= x"CC220008";
end if;
if pc = 7640 then
	inst <= x"022001DC";
end if;
if pc = 7644 then
	inst <= x"C43C0030";
end if;
if pc = 7648 then
	inst <= x"C17DFFFC";
end if;
if pc = 7652 then
	inst <= x"03DC003C";
end if;
if pc = 7656 then
	inst <= x"037E000C";
end if;
if pc = 7660 then
	inst <= x"C57DFFFC";
end if;
if pc = 7664 then
	inst <= x"820007C0";
end if;
if pc = 7668 then
	inst <= x"07DC003C";
end if;
if pc = 7672 then
	inst <= x"C03C0030";
end if;
if pc = 7676 then
	inst <= x"CC220000";
end if;
if pc = 7680 then
	inst <= x"C1FDFFFC";
end if;
if pc = 7684 then
	inst <= x"C8240000";
end if;
if pc = 7688 then
	inst <= x"C8400098";
end if;
if pc = 7692 then
	inst <= x"C43C0000";
end if;
if pc = 7696 then
	inst <= x"CC5C0008";
end if;
if pc = 7700 then
	inst <= x"C45C0010";
end if;
if pc = 7704 then
	inst <= x"8E241E3C";
end if;
if pc = 7708 then
	inst <= x"44224000";
end if;
if pc = 7712 then
	inst <= x"C17DFFFC";
end if;
if pc = 7716 then
	inst <= x"03DC001C";
end if;
if pc = 7720 then
	inst <= x"037E000C";
end if;
if pc = 7724 then
	inst <= x"C57DFFFC";
end if;
if pc = 7728 then
	inst <= x"82001270";
end if;
if pc = 7732 then
	inst <= x"07DC001C";
end if;
if pc = 7736 then
	inst <= x"82001EAC";
end if;
if pc = 7740 then
	inst <= x"8E021E8C";
end if;
if pc = 7744 then
	inst <= x"C8600090";
end if;
if pc = 7748 then
	inst <= x"8E621E68";
end if;
if pc = 7752 then
	inst <= x"40224000";
end if;
if pc = 7756 then
	inst <= x"C17DFFFC";
end if;
if pc = 7760 then
	inst <= x"03DC001C";
end if;
if pc = 7764 then
	inst <= x"037E000C";
end if;
if pc = 7768 then
	inst <= x"C57DFFFC";
end if;
if pc = 7772 then
	inst <= x"82001270";
end if;
if pc = 7776 then
	inst <= x"07DC001C";
end if;
if pc = 7780 then
	inst <= x"82001E88";
end if;
if pc = 7784 then
	inst <= x"02600001";
end if;
if pc = 7788 then
	inst <= x"C17DFFFC";
end if;
if pc = 7792 then
	inst <= x"00260000";
end if;
if pc = 7796 then
	inst <= x"03DC001C";
end if;
if pc = 7800 then
	inst <= x"037E000C";
end if;
if pc = 7804 then
	inst <= x"C57DFFFC";
end if;
if pc = 7808 then
	inst <= x"82000B88";
end if;
if pc = 7812 then
	inst <= x"07DC001C";
end if;
if pc = 7816 then
	inst <= x"82001EAC";
end if;
if pc = 7820 then
	inst <= x"0260FFFF";
end if;
if pc = 7824 then
	inst <= x"C17DFFFC";
end if;
if pc = 7828 then
	inst <= x"00260000";
end if;
if pc = 7832 then
	inst <= x"03DC001C";
end if;
if pc = 7836 then
	inst <= x"037E000C";
end if;
if pc = 7840 then
	inst <= x"C57DFFFC";
end if;
if pc = 7844 then
	inst <= x"82000B88";
end if;
if pc = 7848 then
	inst <= x"07DC001C";
end if;
if pc = 7852 then
	inst <= x"C03C0010";
end if;
if pc = 7856 then
	inst <= x"C8420000";
end if;
if pc = 7860 then
	inst <= x"C87C0008";
end if;
if pc = 7864 then
	inst <= x"CC3C0018";
end if;
if pc = 7868 then
	inst <= x"8E461EE4";
end if;
if pc = 7872 then
	inst <= x"44446000";
end if;
if pc = 7876 then
	inst <= x"C17DFFFC";
end if;
if pc = 7880 then
	inst <= x"40204000";
end if;
if pc = 7884 then
	inst <= x"03DC0028";
end if;
if pc = 7888 then
	inst <= x"037E000C";
end if;
if pc = 7892 then
	inst <= x"C57DFFFC";
end if;
if pc = 7896 then
	inst <= x"82000EC4";
end if;
if pc = 7900 then
	inst <= x"07DC0028";
end if;
if pc = 7904 then
	inst <= x"82001F60";
end if;
if pc = 7908 then
	inst <= x"8E041F3C";
end if;
if pc = 7912 then
	inst <= x"C8800090";
end if;
if pc = 7916 then
	inst <= x"8E841F14";
end if;
if pc = 7920 then
	inst <= x"40446000";
end if;
if pc = 7924 then
	inst <= x"C17DFFFC";
end if;
if pc = 7928 then
	inst <= x"40204000";
end if;
if pc = 7932 then
	inst <= x"03DC0028";
end if;
if pc = 7936 then
	inst <= x"037E000C";
end if;
if pc = 7940 then
	inst <= x"C57DFFFC";
end if;
if pc = 7944 then
	inst <= x"82000EC4";
end if;
if pc = 7948 then
	inst <= x"07DC0028";
end if;
if pc = 7952 then
	inst <= x"82001F38";
end if;
if pc = 7956 then
	inst <= x"02400001";
end if;
if pc = 7960 then
	inst <= x"C17DFFFC";
end if;
if pc = 7964 then
	inst <= x"00240000";
end if;
if pc = 7968 then
	inst <= x"40204000";
end if;
if pc = 7972 then
	inst <= x"03DC0028";
end if;
if pc = 7976 then
	inst <= x"037E000C";
end if;
if pc = 7980 then
	inst <= x"C57DFFFC";
end if;
if pc = 7984 then
	inst <= x"8200084C";
end if;
if pc = 7988 then
	inst <= x"07DC0028";
end if;
if pc = 7992 then
	inst <= x"82001F60";
end if;
if pc = 7996 then
	inst <= x"0240FFFF";
end if;
if pc = 8000 then
	inst <= x"C17DFFFC";
end if;
if pc = 8004 then
	inst <= x"00240000";
end if;
if pc = 8008 then
	inst <= x"40204000";
end if;
if pc = 8012 then
	inst <= x"03DC0028";
end if;
if pc = 8016 then
	inst <= x"037E000C";
end if;
if pc = 8020 then
	inst <= x"C57DFFFC";
end if;
if pc = 8024 then
	inst <= x"8200084C";
end if;
if pc = 8028 then
	inst <= x"07DC0028";
end if;
if pc = 8032 then
	inst <= x"C03C0010";
end if;
if pc = 8036 then
	inst <= x"C8420004";
end if;
if pc = 8040 then
	inst <= x"C87C0008";
end if;
if pc = 8044 then
	inst <= x"CC3C0020";
end if;
if pc = 8048 then
	inst <= x"8E461F98";
end if;
if pc = 8052 then
	inst <= x"44446000";
end if;
if pc = 8056 then
	inst <= x"C17DFFFC";
end if;
if pc = 8060 then
	inst <= x"40204000";
end if;
if pc = 8064 then
	inst <= x"03DC0030";
end if;
if pc = 8068 then
	inst <= x"037E000C";
end if;
if pc = 8072 then
	inst <= x"C57DFFFC";
end if;
if pc = 8076 then
	inst <= x"82001270";
end if;
if pc = 8080 then
	inst <= x"07DC0030";
end if;
if pc = 8084 then
	inst <= x"82002014";
end if;
if pc = 8088 then
	inst <= x"8E041FF0";
end if;
if pc = 8092 then
	inst <= x"C8800090";
end if;
if pc = 8096 then
	inst <= x"8E841FC8";
end if;
if pc = 8100 then
	inst <= x"40446000";
end if;
if pc = 8104 then
	inst <= x"C17DFFFC";
end if;
if pc = 8108 then
	inst <= x"40204000";
end if;
if pc = 8112 then
	inst <= x"03DC0030";
end if;
if pc = 8116 then
	inst <= x"037E000C";
end if;
if pc = 8120 then
	inst <= x"C57DFFFC";
end if;
if pc = 8124 then
	inst <= x"82001270";
end if;
if pc = 8128 then
	inst <= x"07DC0030";
end if;
if pc = 8132 then
	inst <= x"82001FEC";
end if;
if pc = 8136 then
	inst <= x"02400001";
end if;
if pc = 8140 then
	inst <= x"C17DFFFC";
end if;
if pc = 8144 then
	inst <= x"00240000";
end if;
if pc = 8148 then
	inst <= x"40204000";
end if;
if pc = 8152 then
	inst <= x"03DC0030";
end if;
if pc = 8156 then
	inst <= x"037E000C";
end if;
if pc = 8160 then
	inst <= x"C57DFFFC";
end if;
if pc = 8164 then
	inst <= x"82000B88";
end if;
if pc = 8168 then
	inst <= x"07DC0030";
end if;
if pc = 8172 then
	inst <= x"82002014";
end if;
if pc = 8176 then
	inst <= x"0240FFFF";
end if;
if pc = 8180 then
	inst <= x"C17DFFFC";
end if;
if pc = 8184 then
	inst <= x"00240000";
end if;
if pc = 8188 then
	inst <= x"40204000";
end if;
if pc = 8192 then
	inst <= x"03DC0030";
end if;
if pc = 8196 then
	inst <= x"037E000C";
end if;
if pc = 8200 then
	inst <= x"C57DFFFC";
end if;
if pc = 8204 then
	inst <= x"82000B88";
end if;
if pc = 8208 then
	inst <= x"07DC0030";
end if;
if pc = 8212 then
	inst <= x"C03C0010";
end if;
if pc = 8216 then
	inst <= x"C8420004";
end if;
if pc = 8220 then
	inst <= x"C87C0008";
end if;
if pc = 8224 then
	inst <= x"CC3C0028";
end if;
if pc = 8228 then
	inst <= x"8E46204C";
end if;
if pc = 8232 then
	inst <= x"44446000";
end if;
if pc = 8236 then
	inst <= x"C17DFFFC";
end if;
if pc = 8240 then
	inst <= x"40204000";
end if;
if pc = 8244 then
	inst <= x"03DC0038";
end if;
if pc = 8248 then
	inst <= x"037E000C";
end if;
if pc = 8252 then
	inst <= x"C57DFFFC";
end if;
if pc = 8256 then
	inst <= x"82000EC4";
end if;
if pc = 8260 then
	inst <= x"07DC0038";
end if;
if pc = 8264 then
	inst <= x"820020C8";
end if;
if pc = 8268 then
	inst <= x"8E0420A4";
end if;
if pc = 8272 then
	inst <= x"C8800090";
end if;
if pc = 8276 then
	inst <= x"8E84207C";
end if;
if pc = 8280 then
	inst <= x"40446000";
end if;
if pc = 8284 then
	inst <= x"C17DFFFC";
end if;
if pc = 8288 then
	inst <= x"40204000";
end if;
if pc = 8292 then
	inst <= x"03DC0038";
end if;
if pc = 8296 then
	inst <= x"037E000C";
end if;
if pc = 8300 then
	inst <= x"C57DFFFC";
end if;
if pc = 8304 then
	inst <= x"82000EC4";
end if;
if pc = 8308 then
	inst <= x"07DC0038";
end if;
if pc = 8312 then
	inst <= x"820020A0";
end if;
if pc = 8316 then
	inst <= x"02400001";
end if;
if pc = 8320 then
	inst <= x"C17DFFFC";
end if;
if pc = 8324 then
	inst <= x"00240000";
end if;
if pc = 8328 then
	inst <= x"40204000";
end if;
if pc = 8332 then
	inst <= x"03DC0038";
end if;
if pc = 8336 then
	inst <= x"037E000C";
end if;
if pc = 8340 then
	inst <= x"C57DFFFC";
end if;
if pc = 8344 then
	inst <= x"8200084C";
end if;
if pc = 8348 then
	inst <= x"07DC0038";
end if;
if pc = 8352 then
	inst <= x"820020C8";
end if;
if pc = 8356 then
	inst <= x"0240FFFF";
end if;
if pc = 8360 then
	inst <= x"C17DFFFC";
end if;
if pc = 8364 then
	inst <= x"00240000";
end if;
if pc = 8368 then
	inst <= x"40204000";
end if;
if pc = 8372 then
	inst <= x"03DC0038";
end if;
if pc = 8376 then
	inst <= x"037E000C";
end if;
if pc = 8380 then
	inst <= x"C57DFFFC";
end if;
if pc = 8384 then
	inst <= x"8200084C";
end if;
if pc = 8388 then
	inst <= x"07DC0038";
end if;
if pc = 8392 then
	inst <= x"C03C0010";
end if;
if pc = 8396 then
	inst <= x"C8420008";
end if;
if pc = 8400 then
	inst <= x"C87C0008";
end if;
if pc = 8404 then
	inst <= x"CC3C0030";
end if;
if pc = 8408 then
	inst <= x"8E462100";
end if;
if pc = 8412 then
	inst <= x"44446000";
end if;
if pc = 8416 then
	inst <= x"C17DFFFC";
end if;
if pc = 8420 then
	inst <= x"40204000";
end if;
if pc = 8424 then
	inst <= x"03DC0040";
end if;
if pc = 8428 then
	inst <= x"037E000C";
end if;
if pc = 8432 then
	inst <= x"C57DFFFC";
end if;
if pc = 8436 then
	inst <= x"82001270";
end if;
if pc = 8440 then
	inst <= x"07DC0040";
end if;
if pc = 8444 then
	inst <= x"8200217C";
end if;
if pc = 8448 then
	inst <= x"8E042158";
end if;
if pc = 8452 then
	inst <= x"C8800090";
end if;
if pc = 8456 then
	inst <= x"8E842130";
end if;
if pc = 8460 then
	inst <= x"40446000";
end if;
if pc = 8464 then
	inst <= x"C17DFFFC";
end if;
if pc = 8468 then
	inst <= x"40204000";
end if;
if pc = 8472 then
	inst <= x"03DC0040";
end if;
if pc = 8476 then
	inst <= x"037E000C";
end if;
if pc = 8480 then
	inst <= x"C57DFFFC";
end if;
if pc = 8484 then
	inst <= x"82001270";
end if;
if pc = 8488 then
	inst <= x"07DC0040";
end if;
if pc = 8492 then
	inst <= x"82002154";
end if;
if pc = 8496 then
	inst <= x"02400001";
end if;
if pc = 8500 then
	inst <= x"C17DFFFC";
end if;
if pc = 8504 then
	inst <= x"00240000";
end if;
if pc = 8508 then
	inst <= x"40204000";
end if;
if pc = 8512 then
	inst <= x"03DC0040";
end if;
if pc = 8516 then
	inst <= x"037E000C";
end if;
if pc = 8520 then
	inst <= x"C57DFFFC";
end if;
if pc = 8524 then
	inst <= x"82000B88";
end if;
if pc = 8528 then
	inst <= x"07DC0040";
end if;
if pc = 8532 then
	inst <= x"8200217C";
end if;
if pc = 8536 then
	inst <= x"0240FFFF";
end if;
if pc = 8540 then
	inst <= x"C17DFFFC";
end if;
if pc = 8544 then
	inst <= x"00240000";
end if;
if pc = 8548 then
	inst <= x"40204000";
end if;
if pc = 8552 then
	inst <= x"03DC0040";
end if;
if pc = 8556 then
	inst <= x"037E000C";
end if;
if pc = 8560 then
	inst <= x"C57DFFFC";
end if;
if pc = 8564 then
	inst <= x"82000B88";
end if;
if pc = 8568 then
	inst <= x"07DC0040";
end if;
if pc = 8572 then
	inst <= x"C03C0010";
end if;
if pc = 8576 then
	inst <= x"C8420008";
end if;
if pc = 8580 then
	inst <= x"C87C0008";
end if;
if pc = 8584 then
	inst <= x"CC3C0038";
end if;
if pc = 8588 then
	inst <= x"8E4621B4";
end if;
if pc = 8592 then
	inst <= x"44446000";
end if;
if pc = 8596 then
	inst <= x"C17DFFFC";
end if;
if pc = 8600 then
	inst <= x"40204000";
end if;
if pc = 8604 then
	inst <= x"03DC0048";
end if;
if pc = 8608 then
	inst <= x"037E000C";
end if;
if pc = 8612 then
	inst <= x"C57DFFFC";
end if;
if pc = 8616 then
	inst <= x"82000EC4";
end if;
if pc = 8620 then
	inst <= x"07DC0048";
end if;
if pc = 8624 then
	inst <= x"82002230";
end if;
if pc = 8628 then
	inst <= x"8E04220C";
end if;
if pc = 8632 then
	inst <= x"C8800090";
end if;
if pc = 8636 then
	inst <= x"8E8421E4";
end if;
if pc = 8640 then
	inst <= x"40446000";
end if;
if pc = 8644 then
	inst <= x"C17DFFFC";
end if;
if pc = 8648 then
	inst <= x"40204000";
end if;
if pc = 8652 then
	inst <= x"03DC0048";
end if;
if pc = 8656 then
	inst <= x"037E000C";
end if;
if pc = 8660 then
	inst <= x"C57DFFFC";
end if;
if pc = 8664 then
	inst <= x"82000EC4";
end if;
if pc = 8668 then
	inst <= x"07DC0048";
end if;
if pc = 8672 then
	inst <= x"82002208";
end if;
if pc = 8676 then
	inst <= x"02400001";
end if;
if pc = 8680 then
	inst <= x"C17DFFFC";
end if;
if pc = 8684 then
	inst <= x"00240000";
end if;
if pc = 8688 then
	inst <= x"40204000";
end if;
if pc = 8692 then
	inst <= x"03DC0048";
end if;
if pc = 8696 then
	inst <= x"037E000C";
end if;
if pc = 8700 then
	inst <= x"C57DFFFC";
end if;
if pc = 8704 then
	inst <= x"8200084C";
end if;
if pc = 8708 then
	inst <= x"07DC0048";
end if;
if pc = 8712 then
	inst <= x"82002230";
end if;
if pc = 8716 then
	inst <= x"0240FFFF";
end if;
if pc = 8720 then
	inst <= x"C17DFFFC";
end if;
if pc = 8724 then
	inst <= x"00240000";
end if;
if pc = 8728 then
	inst <= x"40204000";
end if;
if pc = 8732 then
	inst <= x"03DC0048";
end if;
if pc = 8736 then
	inst <= x"037E000C";
end if;
if pc = 8740 then
	inst <= x"C57DFFFC";
end if;
if pc = 8744 then
	inst <= x"8200084C";
end if;
if pc = 8748 then
	inst <= x"07DC0048";
end if;
if pc = 8752 then
	inst <= x"C85C0038";
end if;
if pc = 8756 then
	inst <= x"C87C0028";
end if;
if pc = 8760 then
	inst <= x"48864000";
end if;
if pc = 8764 then
	inst <= x"C8BC0030";
end if;
if pc = 8768 then
	inst <= x"C8DC0020";
end if;
if pc = 8772 then
	inst <= x"48ECA000";
end if;
if pc = 8776 then
	inst <= x"490E4000";
end if;
if pc = 8780 then
	inst <= x"C93C0018";
end if;
if pc = 8784 then
	inst <= x"49522000";
end if;
if pc = 8788 then
	inst <= x"45114000";
end if;
if pc = 8792 then
	inst <= x"4952A000";
end if;
if pc = 8796 then
	inst <= x"49744000";
end if;
if pc = 8800 then
	inst <= x"498C2000";
end if;
if pc = 8804 then
	inst <= x"41778000";
end if;
if pc = 8808 then
	inst <= x"49862000";
end if;
if pc = 8812 then
	inst <= x"48EE2000";
end if;
if pc = 8816 then
	inst <= x"49B24000";
end if;
if pc = 8820 then
	inst <= x"40EFA000";
end if;
if pc = 8824 then
	inst <= x"48342000";
end if;
if pc = 8828 then
	inst <= x"484C4000";
end if;
if pc = 8832 then
	inst <= x"44224000";
end if;
if pc = 8836 then
	inst <= x"4440A000";
end if;
if pc = 8840 then
	inst <= x"48AC6000";
end if;
if pc = 8844 then
	inst <= x"48726000";
end if;
if pc = 8848 then
	inst <= x"C03C0000";
end if;
if pc = 8852 then
	inst <= x"C8C20000";
end if;
if pc = 8856 then
	inst <= x"C9220004";
end if;
if pc = 8860 then
	inst <= x"C9420008";
end if;
if pc = 8864 then
	inst <= x"49A88000";
end if;
if pc = 8868 then
	inst <= x"49ADA000";
end if;
if pc = 8872 then
	inst <= x"49D98000";
end if;
if pc = 8876 then
	inst <= x"49D3C000";
end if;
if pc = 8880 then
	inst <= x"41BBC000";
end if;
if pc = 8884 then
	inst <= x"49C44000";
end if;
if pc = 8888 then
	inst <= x"49D5C000";
end if;
if pc = 8892 then
	inst <= x"41BBC000";
end if;
if pc = 8896 then
	inst <= x"CDA20000";
end if;
if pc = 8900 then
	inst <= x"49B10000";
end if;
if pc = 8904 then
	inst <= x"49ADA000";
end if;
if pc = 8908 then
	inst <= x"49CEE000";
end if;
if pc = 8912 then
	inst <= x"49D3C000";
end if;
if pc = 8916 then
	inst <= x"41BBC000";
end if;
if pc = 8920 then
	inst <= x"49CAA000";
end if;
if pc = 8924 then
	inst <= x"49D5C000";
end if;
if pc = 8928 then
	inst <= x"41BBC000";
end if;
if pc = 8932 then
	inst <= x"CDA20004";
end if;
if pc = 8936 then
	inst <= x"49B76000";
end if;
if pc = 8940 then
	inst <= x"49ADA000";
end if;
if pc = 8944 then
	inst <= x"49C22000";
end if;
if pc = 8948 then
	inst <= x"49D3C000";
end if;
if pc = 8952 then
	inst <= x"41BBC000";
end if;
if pc = 8956 then
	inst <= x"49C66000";
end if;
if pc = 8960 then
	inst <= x"49D5C000";
end if;
if pc = 8964 then
	inst <= x"41BBC000";
end if;
if pc = 8968 then
	inst <= x"CDA20008";
end if;
if pc = 8972 then
	inst <= x"C9A00080";
end if;
if pc = 8976 then
	inst <= x"49CD0000";
end if;
if pc = 8980 then
	inst <= x"49DD6000";
end if;
if pc = 8984 then
	inst <= x"49F2E000";
end if;
if pc = 8988 then
	inst <= x"49FE2000";
end if;
if pc = 8992 then
	inst <= x"41DDE000";
end if;
if pc = 8996 then
	inst <= x"49F4A000";
end if;
if pc = 9000 then
	inst <= x"49FE6000";
end if;
if pc = 9004 then
	inst <= x"41DDE000";
end if;
if pc = 9008 then
	inst <= x"49DBC000";
end if;
if pc = 9012 then
	inst <= x"C03C0010";
end if;
if pc = 9016 then
	inst <= x"CDC20000";
end if;
if pc = 9020 then
	inst <= x"488C8000";
end if;
if pc = 9024 then
	inst <= x"48C96000";
end if;
if pc = 9028 then
	inst <= x"49338000";
end if;
if pc = 9032 then
	inst <= x"48322000";
end if;
if pc = 9036 then
	inst <= x"402C2000";
end if;
if pc = 9040 then
	inst <= x"48544000";
end if;
if pc = 9044 then
	inst <= x"48646000";
end if;
if pc = 9048 then
	inst <= x"40226000";
end if;
if pc = 9052 then
	inst <= x"483A2000";
end if;
if pc = 9056 then
	inst <= x"CC220004";
end if;
if pc = 9060 then
	inst <= x"48290000";
end if;
if pc = 9064 then
	inst <= x"4872E000";
end if;
if pc = 9068 then
	inst <= x"40226000";
end if;
if pc = 9072 then
	inst <= x"4844A000";
end if;
if pc = 9076 then
	inst <= x"40224000";
end if;
if pc = 9080 then
	inst <= x"483A2000";
end if;
if pc = 9084 then
	inst <= x"CC220008";
end if;
if pc = 9088 then
	inst <= x"C1FDFFFC";
end if;
if pc = 9092 then
	inst <= x"C43C0000";
end if;
if pc = 9096 then
	inst <= x"C17DFFFC";
end if;
if pc = 9100 then
	inst <= x"03DC000C";
end if;
if pc = 9104 then
	inst <= x"037E000C";
end if;
if pc = 9108 then
	inst <= x"C57DFFFC";
end if;
if pc = 9112 then
	inst <= x"82000794";
end if;
if pc = 9116 then
	inst <= x"07DC000C";
end if;
if pc = 9120 then
	inst <= x"0240FFFF";
end if;
if pc = 9124 then
	inst <= x"82242928";
end if;
if pc = 9128 then
	inst <= x"C43C0004";
end if;
if pc = 9132 then
	inst <= x"C17DFFFC";
end if;
if pc = 9136 then
	inst <= x"03DC0010";
end if;
if pc = 9140 then
	inst <= x"037E000C";
end if;
if pc = 9144 then
	inst <= x"C57DFFFC";
end if;
if pc = 9148 then
	inst <= x"82000794";
end if;
if pc = 9152 then
	inst <= x"07DC0010";
end if;
if pc = 9156 then
	inst <= x"C43C0008";
end if;
if pc = 9160 then
	inst <= x"C17DFFFC";
end if;
if pc = 9164 then
	inst <= x"03DC0014";
end if;
if pc = 9168 then
	inst <= x"037E000C";
end if;
if pc = 9172 then
	inst <= x"C57DFFFC";
end if;
if pc = 9176 then
	inst <= x"82000794";
end if;
if pc = 9180 then
	inst <= x"07DC0014";
end if;
if pc = 9184 then
	inst <= x"C43C000C";
end if;
if pc = 9188 then
	inst <= x"C17DFFFC";
end if;
if pc = 9192 then
	inst <= x"03DC0018";
end if;
if pc = 9196 then
	inst <= x"037E000C";
end if;
if pc = 9200 then
	inst <= x"C57DFFFC";
end if;
if pc = 9204 then
	inst <= x"82000794";
end if;
if pc = 9208 then
	inst <= x"07DC0018";
end if;
if pc = 9212 then
	inst <= x"02400003";
end if;
if pc = 9216 then
	inst <= x"40200000";
end if;
if pc = 9220 then
	inst <= x"C43C0010";
end if;
if pc = 9224 then
	inst <= x"CC3C0018";
end if;
if pc = 9228 then
	inst <= x"C17DFFFC";
end if;
if pc = 9232 then
	inst <= x"00240000";
end if;
if pc = 9236 then
	inst <= x"03DC0028";
end if;
if pc = 9240 then
	inst <= x"037E000C";
end if;
if pc = 9244 then
	inst <= x"C57DFFFC";
end if;
if pc = 9248 then
	inst <= x"8200081C";
end if;
if pc = 9252 then
	inst <= x"07DC0028";
end if;
if pc = 9256 then
	inst <= x"C43C0020";
end if;
if pc = 9260 then
	inst <= x"C17DFFFC";
end if;
if pc = 9264 then
	inst <= x"03DC002C";
end if;
if pc = 9268 then
	inst <= x"037E000C";
end if;
if pc = 9272 then
	inst <= x"C57DFFFC";
end if;
if pc = 9276 then
	inst <= x"820007C0";
end if;
if pc = 9280 then
	inst <= x"07DC002C";
end if;
if pc = 9284 then
	inst <= x"C03C0020";
end if;
if pc = 9288 then
	inst <= x"CC220000";
end if;
if pc = 9292 then
	inst <= x"C17DFFFC";
end if;
if pc = 9296 then
	inst <= x"03DC002C";
end if;
if pc = 9300 then
	inst <= x"037E000C";
end if;
if pc = 9304 then
	inst <= x"C57DFFFC";
end if;
if pc = 9308 then
	inst <= x"820007C0";
end if;
if pc = 9312 then
	inst <= x"07DC002C";
end if;
if pc = 9316 then
	inst <= x"C03C0020";
end if;
if pc = 9320 then
	inst <= x"CC220004";
end if;
if pc = 9324 then
	inst <= x"C17DFFFC";
end if;
if pc = 9328 then
	inst <= x"03DC002C";
end if;
if pc = 9332 then
	inst <= x"037E000C";
end if;
if pc = 9336 then
	inst <= x"C57DFFFC";
end if;
if pc = 9340 then
	inst <= x"820007C0";
end if;
if pc = 9344 then
	inst <= x"07DC002C";
end if;
if pc = 9348 then
	inst <= x"C03C0020";
end if;
if pc = 9352 then
	inst <= x"CC220008";
end if;
if pc = 9356 then
	inst <= x"02400003";
end if;
if pc = 9360 then
	inst <= x"C83C0018";
end if;
if pc = 9364 then
	inst <= x"C17DFFFC";
end if;
if pc = 9368 then
	inst <= x"00240000";
end if;
if pc = 9372 then
	inst <= x"03DC002C";
end if;
if pc = 9376 then
	inst <= x"037E000C";
end if;
if pc = 9380 then
	inst <= x"C57DFFFC";
end if;
if pc = 9384 then
	inst <= x"8200081C";
end if;
if pc = 9388 then
	inst <= x"07DC002C";
end if;
if pc = 9392 then
	inst <= x"C43C0024";
end if;
if pc = 9396 then
	inst <= x"C17DFFFC";
end if;
if pc = 9400 then
	inst <= x"03DC0030";
end if;
if pc = 9404 then
	inst <= x"037E000C";
end if;
if pc = 9408 then
	inst <= x"C57DFFFC";
end if;
if pc = 9412 then
	inst <= x"820007C0";
end if;
if pc = 9416 then
	inst <= x"07DC0030";
end if;
if pc = 9420 then
	inst <= x"C03C0024";
end if;
if pc = 9424 then
	inst <= x"CC220000";
end if;
if pc = 9428 then
	inst <= x"C17DFFFC";
end if;
if pc = 9432 then
	inst <= x"03DC0030";
end if;
if pc = 9436 then
	inst <= x"037E000C";
end if;
if pc = 9440 then
	inst <= x"C57DFFFC";
end if;
if pc = 9444 then
	inst <= x"820007C0";
end if;
if pc = 9448 then
	inst <= x"07DC0030";
end if;
if pc = 9452 then
	inst <= x"C03C0024";
end if;
if pc = 9456 then
	inst <= x"CC220004";
end if;
if pc = 9460 then
	inst <= x"C17DFFFC";
end if;
if pc = 9464 then
	inst <= x"03DC0030";
end if;
if pc = 9468 then
	inst <= x"037E000C";
end if;
if pc = 9472 then
	inst <= x"C57DFFFC";
end if;
if pc = 9476 then
	inst <= x"820007C0";
end if;
if pc = 9480 then
	inst <= x"07DC0030";
end if;
if pc = 9484 then
	inst <= x"C03C0024";
end if;
if pc = 9488 then
	inst <= x"CC220008";
end if;
if pc = 9492 then
	inst <= x"C17DFFFC";
end if;
if pc = 9496 then
	inst <= x"03DC0030";
end if;
if pc = 9500 then
	inst <= x"037E000C";
end if;
if pc = 9504 then
	inst <= x"C57DFFFC";
end if;
if pc = 9508 then
	inst <= x"820007C0";
end if;
if pc = 9512 then
	inst <= x"07DC0030";
end if;
if pc = 9516 then
	inst <= x"8E202538";
end if;
if pc = 9520 then
	inst <= x"02200000";
end if;
if pc = 9524 then
	inst <= x"8200253C";
end if;
if pc = 9528 then
	inst <= x"02200001";
end if;
if pc = 9532 then
	inst <= x"02400002";
end if;
if pc = 9536 then
	inst <= x"C85C0018";
end if;
if pc = 9540 then
	inst <= x"CC3C0028";
end if;
if pc = 9544 then
	inst <= x"C43C0030";
end if;
if pc = 9548 then
	inst <= x"C17DFFFC";
end if;
if pc = 9552 then
	inst <= x"00240000";
end if;
if pc = 9556 then
	inst <= x"40204000";
end if;
if pc = 9560 then
	inst <= x"03DC003C";
end if;
if pc = 9564 then
	inst <= x"037E000C";
end if;
if pc = 9568 then
	inst <= x"C57DFFFC";
end if;
if pc = 9572 then
	inst <= x"8200081C";
end if;
if pc = 9576 then
	inst <= x"07DC003C";
end if;
if pc = 9580 then
	inst <= x"C43C0034";
end if;
if pc = 9584 then
	inst <= x"C17DFFFC";
end if;
if pc = 9588 then
	inst <= x"03DC0040";
end if;
if pc = 9592 then
	inst <= x"037E000C";
end if;
if pc = 9596 then
	inst <= x"C57DFFFC";
end if;
if pc = 9600 then
	inst <= x"820007C0";
end if;
if pc = 9604 then
	inst <= x"07DC0040";
end if;
if pc = 9608 then
	inst <= x"C03C0034";
end if;
if pc = 9612 then
	inst <= x"CC220000";
end if;
if pc = 9616 then
	inst <= x"C17DFFFC";
end if;
if pc = 9620 then
	inst <= x"03DC0040";
end if;
if pc = 9624 then
	inst <= x"037E000C";
end if;
if pc = 9628 then
	inst <= x"C57DFFFC";
end if;
if pc = 9632 then
	inst <= x"820007C0";
end if;
if pc = 9636 then
	inst <= x"07DC0040";
end if;
if pc = 9640 then
	inst <= x"C03C0034";
end if;
if pc = 9644 then
	inst <= x"CC220004";
end if;
if pc = 9648 then
	inst <= x"02400003";
end if;
if pc = 9652 then
	inst <= x"C83C0018";
end if;
if pc = 9656 then
	inst <= x"C17DFFFC";
end if;
if pc = 9660 then
	inst <= x"00240000";
end if;
if pc = 9664 then
	inst <= x"03DC0040";
end if;
if pc = 9668 then
	inst <= x"037E000C";
end if;
if pc = 9672 then
	inst <= x"C57DFFFC";
end if;
if pc = 9676 then
	inst <= x"8200081C";
end if;
if pc = 9680 then
	inst <= x"07DC0040";
end if;
if pc = 9684 then
	inst <= x"C43C0038";
end if;
if pc = 9688 then
	inst <= x"C17DFFFC";
end if;
if pc = 9692 then
	inst <= x"03DC0044";
end if;
if pc = 9696 then
	inst <= x"037E000C";
end if;
if pc = 9700 then
	inst <= x"C57DFFFC";
end if;
if pc = 9704 then
	inst <= x"820007C0";
end if;
if pc = 9708 then
	inst <= x"07DC0044";
end if;
if pc = 9712 then
	inst <= x"C03C0038";
end if;
if pc = 9716 then
	inst <= x"CC220000";
end if;
if pc = 9720 then
	inst <= x"C17DFFFC";
end if;
if pc = 9724 then
	inst <= x"03DC0044";
end if;
if pc = 9728 then
	inst <= x"037E000C";
end if;
if pc = 9732 then
	inst <= x"C57DFFFC";
end if;
if pc = 9736 then
	inst <= x"820007C0";
end if;
if pc = 9740 then
	inst <= x"07DC0044";
end if;
if pc = 9744 then
	inst <= x"C03C0038";
end if;
if pc = 9748 then
	inst <= x"CC220004";
end if;
if pc = 9752 then
	inst <= x"C17DFFFC";
end if;
if pc = 9756 then
	inst <= x"03DC0044";
end if;
if pc = 9760 then
	inst <= x"037E000C";
end if;
if pc = 9764 then
	inst <= x"C57DFFFC";
end if;
if pc = 9768 then
	inst <= x"820007C0";
end if;
if pc = 9772 then
	inst <= x"07DC0044";
end if;
if pc = 9776 then
	inst <= x"C03C0038";
end if;
if pc = 9780 then
	inst <= x"CC220008";
end if;
if pc = 9784 then
	inst <= x"02400003";
end if;
if pc = 9788 then
	inst <= x"C83C0018";
end if;
if pc = 9792 then
	inst <= x"C17DFFFC";
end if;
if pc = 9796 then
	inst <= x"00240000";
end if;
if pc = 9800 then
	inst <= x"03DC0044";
end if;
if pc = 9804 then
	inst <= x"037E000C";
end if;
if pc = 9808 then
	inst <= x"C57DFFFC";
end if;
if pc = 9812 then
	inst <= x"8200081C";
end if;
if pc = 9816 then
	inst <= x"07DC0044";
end if;
if pc = 9820 then
	inst <= x"C05C0010";
end if;
if pc = 9824 then
	inst <= x"824026E8";
end if;
if pc = 9828 then
	inst <= x"C43C003C";
end if;
if pc = 9832 then
	inst <= x"C17DFFFC";
end if;
if pc = 9836 then
	inst <= x"03DC0048";
end if;
if pc = 9840 then
	inst <= x"037E000C";
end if;
if pc = 9844 then
	inst <= x"C57DFFFC";
end if;
if pc = 9848 then
	inst <= x"820007C0";
end if;
if pc = 9852 then
	inst <= x"07DC0048";
end if;
if pc = 9856 then
	inst <= x"C840008C";
end if;
if pc = 9860 then
	inst <= x"48224000";
end if;
if pc = 9864 then
	inst <= x"C03C003C";
end if;
if pc = 9868 then
	inst <= x"CC220000";
end if;
if pc = 9872 then
	inst <= x"CC5C0040";
end if;
if pc = 9876 then
	inst <= x"C17DFFFC";
end if;
if pc = 9880 then
	inst <= x"03DC0050";
end if;
if pc = 9884 then
	inst <= x"037E000C";
end if;
if pc = 9888 then
	inst <= x"C57DFFFC";
end if;
if pc = 9892 then
	inst <= x"820007C0";
end if;
if pc = 9896 then
	inst <= x"07DC0050";
end if;
if pc = 9900 then
	inst <= x"C85C0040";
end if;
if pc = 9904 then
	inst <= x"48224000";
end if;
if pc = 9908 then
	inst <= x"C03C003C";
end if;
if pc = 9912 then
	inst <= x"CC220004";
end if;
if pc = 9916 then
	inst <= x"C17DFFFC";
end if;
if pc = 9920 then
	inst <= x"03DC0050";
end if;
if pc = 9924 then
	inst <= x"037E000C";
end if;
if pc = 9928 then
	inst <= x"C57DFFFC";
end if;
if pc = 9932 then
	inst <= x"820007C0";
end if;
if pc = 9936 then
	inst <= x"07DC0050";
end if;
if pc = 9940 then
	inst <= x"C85C0040";
end if;
if pc = 9944 then
	inst <= x"48224000";
end if;
if pc = 9948 then
	inst <= x"C03C003C";
end if;
if pc = 9952 then
	inst <= x"CC220008";
end if;
if pc = 9956 then
	inst <= x"820026E8";
end if;
if pc = 9960 then
	inst <= x"02400002";
end if;
if pc = 9964 then
	inst <= x"C07C0008";
end if;
if pc = 9968 then
	inst <= x"826426FC";
end if;
if pc = 9972 then
	inst <= x"C05C0030";
end if;
if pc = 9976 then
	inst <= x"82002700";
end if;
if pc = 9980 then
	inst <= x"02400001";
end if;
if pc = 9984 then
	inst <= x"02800004";
end if;
if pc = 9988 then
	inst <= x"C83C0018";
end if;
if pc = 9992 then
	inst <= x"C45C0048";
end if;
if pc = 9996 then
	inst <= x"C43C003C";
end if;
if pc = 10000 then
	inst <= x"C17DFFFC";
end if;
if pc = 10004 then
	inst <= x"00280000";
end if;
if pc = 10008 then
	inst <= x"03DC0054";
end if;
if pc = 10012 then
	inst <= x"037E000C";
end if;
if pc = 10016 then
	inst <= x"C57DFFFC";
end if;
if pc = 10020 then
	inst <= x"8200081C";
end if;
if pc = 10024 then
	inst <= x"07DC0054";
end if;
if pc = 10028 then
	inst <= x"005A0000";
end if;
if pc = 10032 then
	inst <= x"03BA002C";
end if;
if pc = 10036 then
	inst <= x"C4240028";
end if;
if pc = 10040 then
	inst <= x"C03C003C";
end if;
if pc = 10044 then
	inst <= x"C4240024";
end if;
if pc = 10048 then
	inst <= x"C07C0038";
end if;
if pc = 10052 then
	inst <= x"C4640020";
end if;
if pc = 10056 then
	inst <= x"C07C0034";
end if;
if pc = 10060 then
	inst <= x"C464001C";
end if;
if pc = 10064 then
	inst <= x"C07C0048";
end if;
if pc = 10068 then
	inst <= x"C4640018";
end if;
if pc = 10072 then
	inst <= x"C07C0024";
end if;
if pc = 10076 then
	inst <= x"C4640014";
end if;
if pc = 10080 then
	inst <= x"C07C0020";
end if;
if pc = 10084 then
	inst <= x"C4640010";
end if;
if pc = 10088 then
	inst <= x"C09C0010";
end if;
if pc = 10092 then
	inst <= x"C484000C";
end if;
if pc = 10096 then
	inst <= x"C0BC000C";
end if;
if pc = 10100 then
	inst <= x"C4A40008";
end if;
if pc = 10104 then
	inst <= x"C0BC0008";
end if;
if pc = 10108 then
	inst <= x"C4A40004";
end if;
if pc = 10112 then
	inst <= x"C0DC0004";
end if;
if pc = 10116 then
	inst <= x"C4C40000";
end if;
if pc = 10120 then
	inst <= x"02C000C8";
end if;
if pc = 10124 then
	inst <= x"C0FC0000";
end if;
if pc = 10128 then
	inst <= x"22EE0220";
end if;
if pc = 10132 then
	inst <= x"D44CE000";
end if;
if pc = 10136 then
	inst <= x"02400003";
end if;
if pc = 10140 then
	inst <= x"82A427E0";
end if;
if pc = 10144 then
	inst <= x"02400002";
end if;
if pc = 10148 then
	inst <= x"82A427AC";
end if;
if pc = 10152 then
	inst <= x"820027DC";
end if;
if pc = 10156 then
	inst <= x"C83C0028";
end if;
if pc = 10160 then
	inst <= x"8E2027BC";
end if;
if pc = 10164 then
	inst <= x"02400001";
end if;
if pc = 10168 then
	inst <= x"820027C0";
end if;
if pc = 10172 then
	inst <= x"02400000";
end if;
if pc = 10176 then
	inst <= x"C17DFFFC";
end if;
if pc = 10180 then
	inst <= x"00260000";
end if;
if pc = 10184 then
	inst <= x"03DC0054";
end if;
if pc = 10188 then
	inst <= x"037E000C";
end if;
if pc = 10192 then
	inst <= x"C57DFFFC";
end if;
if pc = 10196 then
	inst <= x"8200161C";
end if;
if pc = 10200 then
	inst <= x"07DC0054";
end if;
if pc = 10204 then
	inst <= x"820028F4";
end if;
if pc = 10208 then
	inst <= x"C8260000";
end if;
if pc = 10212 then
	inst <= x"8A202830";
end if;
if pc = 10216 then
	inst <= x"8A202800";
end if;
if pc = 10220 then
	inst <= x"8E0227F8";
end if;
if pc = 10224 then
	inst <= x"C840007C";
end if;
if pc = 10228 then
	inst <= x"820027FC";
end if;
if pc = 10232 then
	inst <= x"C84000A8";
end if;
if pc = 10236 then
	inst <= x"82002804";
end if;
if pc = 10240 then
	inst <= x"40400000";
end if;
if pc = 10244 then
	inst <= x"48222000";
end if;
if pc = 10248 then
	inst <= x"CC5C0050";
end if;
if pc = 10252 then
	inst <= x"C17DFFFC";
end if;
if pc = 10256 then
	inst <= x"03DC0060";
end if;
if pc = 10260 then
	inst <= x"037E000C";
end if;
if pc = 10264 then
	inst <= x"C57DFFFC";
end if;
if pc = 10268 then
	inst <= x"82000844";
end if;
if pc = 10272 then
	inst <= x"07DC0060";
end if;
if pc = 10276 then
	inst <= x"C85C0050";
end if;
if pc = 10280 then
	inst <= x"48242000";
end if;
if pc = 10284 then
	inst <= x"82002834";
end if;
if pc = 10288 then
	inst <= x"40200000";
end if;
if pc = 10292 then
	inst <= x"C03C0020";
end if;
if pc = 10296 then
	inst <= x"CC220000";
end if;
if pc = 10300 then
	inst <= x"C8220004";
end if;
if pc = 10304 then
	inst <= x"8A20288C";
end if;
if pc = 10308 then
	inst <= x"8A20285C";
end if;
if pc = 10312 then
	inst <= x"8E022854";
end if;
if pc = 10316 then
	inst <= x"C840007C";
end if;
if pc = 10320 then
	inst <= x"82002858";
end if;
if pc = 10324 then
	inst <= x"C84000A8";
end if;
if pc = 10328 then
	inst <= x"82002860";
end if;
if pc = 10332 then
	inst <= x"40400000";
end if;
if pc = 10336 then
	inst <= x"48222000";
end if;
if pc = 10340 then
	inst <= x"CC5C0058";
end if;
if pc = 10344 then
	inst <= x"C17DFFFC";
end if;
if pc = 10348 then
	inst <= x"03DC0068";
end if;
if pc = 10352 then
	inst <= x"037E000C";
end if;
if pc = 10356 then
	inst <= x"C57DFFFC";
end if;
if pc = 10360 then
	inst <= x"82000844";
end if;
if pc = 10364 then
	inst <= x"07DC0068";
end if;
if pc = 10368 then
	inst <= x"C85C0058";
end if;
if pc = 10372 then
	inst <= x"48242000";
end if;
if pc = 10376 then
	inst <= x"82002890";
end if;
if pc = 10380 then
	inst <= x"40200000";
end if;
if pc = 10384 then
	inst <= x"C03C0020";
end if;
if pc = 10388 then
	inst <= x"CC220004";
end if;
if pc = 10392 then
	inst <= x"C8220008";
end if;
if pc = 10396 then
	inst <= x"8A2028E8";
end if;
if pc = 10400 then
	inst <= x"8A2028B8";
end if;
if pc = 10404 then
	inst <= x"8E0228B0";
end if;
if pc = 10408 then
	inst <= x"C840007C";
end if;
if pc = 10412 then
	inst <= x"820028B4";
end if;
if pc = 10416 then
	inst <= x"C84000A8";
end if;
if pc = 10420 then
	inst <= x"820028BC";
end if;
if pc = 10424 then
	inst <= x"40400000";
end if;
if pc = 10428 then
	inst <= x"48222000";
end if;
if pc = 10432 then
	inst <= x"CC5C0060";
end if;
if pc = 10436 then
	inst <= x"C17DFFFC";
end if;
if pc = 10440 then
	inst <= x"03DC0070";
end if;
if pc = 10444 then
	inst <= x"037E000C";
end if;
if pc = 10448 then
	inst <= x"C57DFFFC";
end if;
if pc = 10452 then
	inst <= x"82000844";
end if;
if pc = 10456 then
	inst <= x"07DC0070";
end if;
if pc = 10460 then
	inst <= x"C85C0060";
end if;
if pc = 10464 then
	inst <= x"48242000";
end if;
if pc = 10468 then
	inst <= x"820028EC";
end if;
if pc = 10472 then
	inst <= x"40200000";
end if;
if pc = 10476 then
	inst <= x"C03C0020";
end if;
if pc = 10480 then
	inst <= x"CC220008";
end if;
if pc = 10484 then
	inst <= x"C03C0010";
end if;
if pc = 10488 then
	inst <= x"82202920";
end if;
if pc = 10492 then
	inst <= x"C03C0020";
end if;
if pc = 10496 then
	inst <= x"C05C003C";
end if;
if pc = 10500 then
	inst <= x"C17DFFFC";
end if;
if pc = 10504 then
	inst <= x"03DC0070";
end if;
if pc = 10508 then
	inst <= x"037E000C";
end if;
if pc = 10512 then
	inst <= x"C57DFFFC";
end if;
if pc = 10516 then
	inst <= x"82001E04";
end if;
if pc = 10520 then
	inst <= x"07DC0070";
end if;
if pc = 10524 then
	inst <= x"82002920";
end if;
if pc = 10528 then
	inst <= x"02200001";
end if;
if pc = 10532 then
	inst <= x"C1FDFFFC";
end if;
if pc = 10536 then
	inst <= x"02200000";
end if;
if pc = 10540 then
	inst <= x"C1FDFFFC";
end if;
if pc = 10544 then
	inst <= x"0240003C";
end if;
if pc = 10548 then
	inst <= x"8624293C";
end if;
if pc = 10552 then
	inst <= x"C1FDFFFC";
end if;
if pc = 10556 then
	inst <= x"C43C0000";
end if;
if pc = 10560 then
	inst <= x"C17DFFFC";
end if;
if pc = 10564 then
	inst <= x"03DC000C";
end if;
if pc = 10568 then
	inst <= x"037E000C";
end if;
if pc = 10572 then
	inst <= x"C57DFFFC";
end if;
if pc = 10576 then
	inst <= x"82002384";
end if;
if pc = 10580 then
	inst <= x"07DC000C";
end if;
if pc = 10584 then
	inst <= x"82202A34";
end if;
if pc = 10588 then
	inst <= x"C03C0000";
end if;
if pc = 10592 then
	inst <= x"02220001";
end if;
if pc = 10596 then
	inst <= x"0240003C";
end if;
if pc = 10600 then
	inst <= x"86242970";
end if;
if pc = 10604 then
	inst <= x"C1FDFFFC";
end if;
if pc = 10608 then
	inst <= x"C43C0004";
end if;
if pc = 10612 then
	inst <= x"C17DFFFC";
end if;
if pc = 10616 then
	inst <= x"03DC0010";
end if;
if pc = 10620 then
	inst <= x"037E000C";
end if;
if pc = 10624 then
	inst <= x"C57DFFFC";
end if;
if pc = 10628 then
	inst <= x"82002384";
end if;
if pc = 10632 then
	inst <= x"07DC0010";
end if;
if pc = 10636 then
	inst <= x"82202A24";
end if;
if pc = 10640 then
	inst <= x"C03C0004";
end if;
if pc = 10644 then
	inst <= x"02220001";
end if;
if pc = 10648 then
	inst <= x"0240003C";
end if;
if pc = 10652 then
	inst <= x"862429A4";
end if;
if pc = 10656 then
	inst <= x"C1FDFFFC";
end if;
if pc = 10660 then
	inst <= x"C43C0008";
end if;
if pc = 10664 then
	inst <= x"C17DFFFC";
end if;
if pc = 10668 then
	inst <= x"03DC0014";
end if;
if pc = 10672 then
	inst <= x"037E000C";
end if;
if pc = 10676 then
	inst <= x"C57DFFFC";
end if;
if pc = 10680 then
	inst <= x"82002384";
end if;
if pc = 10684 then
	inst <= x"07DC0014";
end if;
if pc = 10688 then
	inst <= x"82202A14";
end if;
if pc = 10692 then
	inst <= x"C03C0008";
end if;
if pc = 10696 then
	inst <= x"02220001";
end if;
if pc = 10700 then
	inst <= x"0240003C";
end if;
if pc = 10704 then
	inst <= x"862429D8";
end if;
if pc = 10708 then
	inst <= x"C1FDFFFC";
end if;
if pc = 10712 then
	inst <= x"C43C000C";
end if;
if pc = 10716 then
	inst <= x"C17DFFFC";
end if;
if pc = 10720 then
	inst <= x"03DC0018";
end if;
if pc = 10724 then
	inst <= x"037E000C";
end if;
if pc = 10728 then
	inst <= x"C57DFFFC";
end if;
if pc = 10732 then
	inst <= x"82002384";
end if;
if pc = 10736 then
	inst <= x"07DC0018";
end if;
if pc = 10740 then
	inst <= x"82202A04";
end if;
if pc = 10744 then
	inst <= x"C03C000C";
end if;
if pc = 10748 then
	inst <= x"02220001";
end if;
if pc = 10752 then
	inst <= x"82002930";
end if;
if pc = 10756 then
	inst <= x"022000C4";
end if;
if pc = 10760 then
	inst <= x"C05C000C";
end if;
if pc = 10764 then
	inst <= x"C4420000";
end if;
if pc = 10768 then
	inst <= x"C1FDFFFC";
end if;
if pc = 10772 then
	inst <= x"022000C4";
end if;
if pc = 10776 then
	inst <= x"C05C0008";
end if;
if pc = 10780 then
	inst <= x"C4420000";
end if;
if pc = 10784 then
	inst <= x"C1FDFFFC";
end if;
if pc = 10788 then
	inst <= x"022000C4";
end if;
if pc = 10792 then
	inst <= x"C05C0004";
end if;
if pc = 10796 then
	inst <= x"C4420000";
end if;
if pc = 10800 then
	inst <= x"C1FDFFFC";
end if;
if pc = 10804 then
	inst <= x"022000C4";
end if;
if pc = 10808 then
	inst <= x"C05C0000";
end if;
if pc = 10812 then
	inst <= x"C4420000";
end if;
if pc = 10816 then
	inst <= x"C1FDFFFC";
end if;
if pc = 10820 then
	inst <= x"C43C0000";
end if;
if pc = 10824 then
	inst <= x"C17DFFFC";
end if;
if pc = 10828 then
	inst <= x"03DC000C";
end if;
if pc = 10832 then
	inst <= x"037E000C";
end if;
if pc = 10836 then
	inst <= x"C57DFFFC";
end if;
if pc = 10840 then
	inst <= x"82000794";
end if;
if pc = 10844 then
	inst <= x"07DC000C";
end if;
if pc = 10848 then
	inst <= x"0240FFFF";
end if;
if pc = 10852 then
	inst <= x"82242BDC";
end if;
if pc = 10856 then
	inst <= x"C05C0000";
end if;
if pc = 10860 then
	inst <= x"02640001";
end if;
if pc = 10864 then
	inst <= x"C43C0004";
end if;
if pc = 10868 then
	inst <= x"C47C0008";
end if;
if pc = 10872 then
	inst <= x"C17DFFFC";
end if;
if pc = 10876 then
	inst <= x"03DC0014";
end if;
if pc = 10880 then
	inst <= x"037E000C";
end if;
if pc = 10884 then
	inst <= x"C57DFFFC";
end if;
if pc = 10888 then
	inst <= x"82000794";
end if;
if pc = 10892 then
	inst <= x"07DC0014";
end if;
if pc = 10896 then
	inst <= x"0240FFFF";
end if;
if pc = 10900 then
	inst <= x"82242BA4";
end if;
if pc = 10904 then
	inst <= x"C05C0008";
end if;
if pc = 10908 then
	inst <= x"02640001";
end if;
if pc = 10912 then
	inst <= x"C43C000C";
end if;
if pc = 10916 then
	inst <= x"C47C0010";
end if;
if pc = 10920 then
	inst <= x"C17DFFFC";
end if;
if pc = 10924 then
	inst <= x"03DC001C";
end if;
if pc = 10928 then
	inst <= x"037E000C";
end if;
if pc = 10932 then
	inst <= x"C57DFFFC";
end if;
if pc = 10936 then
	inst <= x"82000794";
end if;
if pc = 10940 then
	inst <= x"07DC001C";
end if;
if pc = 10944 then
	inst <= x"0240FFFF";
end if;
if pc = 10948 then
	inst <= x"82242B6C";
end if;
if pc = 10952 then
	inst <= x"C05C0010";
end if;
if pc = 10956 then
	inst <= x"02640001";
end if;
if pc = 10960 then
	inst <= x"C43C0014";
end if;
if pc = 10964 then
	inst <= x"C47C0018";
end if;
if pc = 10968 then
	inst <= x"C17DFFFC";
end if;
if pc = 10972 then
	inst <= x"03DC0024";
end if;
if pc = 10976 then
	inst <= x"037E000C";
end if;
if pc = 10980 then
	inst <= x"C57DFFFC";
end if;
if pc = 10984 then
	inst <= x"82000794";
end if;
if pc = 10988 then
	inst <= x"07DC0024";
end if;
if pc = 10992 then
	inst <= x"0240FFFF";
end if;
if pc = 10996 then
	inst <= x"82242B34";
end if;
if pc = 11000 then
	inst <= x"C05C0018";
end if;
if pc = 11004 then
	inst <= x"02640001";
end if;
if pc = 11008 then
	inst <= x"C43C001C";
end if;
if pc = 11012 then
	inst <= x"C17DFFFC";
end if;
if pc = 11016 then
	inst <= x"00260000";
end if;
if pc = 11020 then
	inst <= x"03DC0028";
end if;
if pc = 11024 then
	inst <= x"037E000C";
end if;
if pc = 11028 then
	inst <= x"C57DFFFC";
end if;
if pc = 11032 then
	inst <= x"82002A44";
end if;
if pc = 11036 then
	inst <= x"07DC0028";
end if;
if pc = 11040 then
	inst <= x"C05C0018";
end if;
if pc = 11044 then
	inst <= x"22440220";
end if;
if pc = 11048 then
	inst <= x"C07C001C";
end if;
if pc = 11052 then
	inst <= x"D4624000";
end if;
if pc = 11056 then
	inst <= x"82002B58";
end if;
if pc = 11060 then
	inst <= x"C03C0018";
end if;
if pc = 11064 then
	inst <= x"02220001";
end if;
if pc = 11068 then
	inst <= x"0240FFFF";
end if;
if pc = 11072 then
	inst <= x"C17DFFFC";
end if;
if pc = 11076 then
	inst <= x"03DC0028";
end if;
if pc = 11080 then
	inst <= x"037E000C";
end if;
if pc = 11084 then
	inst <= x"C57DFFFC";
end if;
if pc = 11088 then
	inst <= x"8200081C";
end if;
if pc = 11092 then
	inst <= x"07DC0028";
end if;
if pc = 11096 then
	inst <= x"C05C0010";
end if;
if pc = 11100 then
	inst <= x"22440220";
end if;
if pc = 11104 then
	inst <= x"C07C0014";
end if;
if pc = 11108 then
	inst <= x"D4624000";
end if;
if pc = 11112 then
	inst <= x"82002B90";
end if;
if pc = 11116 then
	inst <= x"C03C0010";
end if;
if pc = 11120 then
	inst <= x"02220001";
end if;
if pc = 11124 then
	inst <= x"0240FFFF";
end if;
if pc = 11128 then
	inst <= x"C17DFFFC";
end if;
if pc = 11132 then
	inst <= x"03DC0028";
end if;
if pc = 11136 then
	inst <= x"037E000C";
end if;
if pc = 11140 then
	inst <= x"C57DFFFC";
end if;
if pc = 11144 then
	inst <= x"8200081C";
end if;
if pc = 11148 then
	inst <= x"07DC0028";
end if;
if pc = 11152 then
	inst <= x"C05C0008";
end if;
if pc = 11156 then
	inst <= x"22440220";
end if;
if pc = 11160 then
	inst <= x"C07C000C";
end if;
if pc = 11164 then
	inst <= x"D4624000";
end if;
if pc = 11168 then
	inst <= x"82002BC8";
end if;
if pc = 11172 then
	inst <= x"C03C0008";
end if;
if pc = 11176 then
	inst <= x"02220001";
end if;
if pc = 11180 then
	inst <= x"0240FFFF";
end if;
if pc = 11184 then
	inst <= x"C17DFFFC";
end if;
if pc = 11188 then
	inst <= x"03DC0028";
end if;
if pc = 11192 then
	inst <= x"037E000C";
end if;
if pc = 11196 then
	inst <= x"C57DFFFC";
end if;
if pc = 11200 then
	inst <= x"8200081C";
end if;
if pc = 11204 then
	inst <= x"07DC0028";
end if;
if pc = 11208 then
	inst <= x"C05C0000";
end if;
if pc = 11212 then
	inst <= x"22440220";
end if;
if pc = 11216 then
	inst <= x"C07C0004";
end if;
if pc = 11220 then
	inst <= x"D4624000";
end if;
if pc = 11224 then
	inst <= x"C1FDFFFC";
end if;
if pc = 11228 then
	inst <= x"C03C0000";
end if;
if pc = 11232 then
	inst <= x"02220001";
end if;
if pc = 11236 then
	inst <= x"0240FFFF";
end if;
if pc = 11240 then
	inst <= x"8200081C";
end if;
if pc = 11244 then
	inst <= x"C43C0000";
end if;
if pc = 11248 then
	inst <= x"C17DFFFC";
end if;
if pc = 11252 then
	inst <= x"03DC000C";
end if;
if pc = 11256 then
	inst <= x"037E000C";
end if;
if pc = 11260 then
	inst <= x"C57DFFFC";
end if;
if pc = 11264 then
	inst <= x"82000794";
end if;
if pc = 11268 then
	inst <= x"07DC000C";
end if;
if pc = 11272 then
	inst <= x"0240FFFF";
end if;
if pc = 11276 then
	inst <= x"82242CE4";
end if;
if pc = 11280 then
	inst <= x"C43C0004";
end if;
if pc = 11284 then
	inst <= x"C17DFFFC";
end if;
if pc = 11288 then
	inst <= x"03DC0010";
end if;
if pc = 11292 then
	inst <= x"037E000C";
end if;
if pc = 11296 then
	inst <= x"C57DFFFC";
end if;
if pc = 11300 then
	inst <= x"82000794";
end if;
if pc = 11304 then
	inst <= x"07DC0010";
end if;
if pc = 11308 then
	inst <= x"0240FFFF";
end if;
if pc = 11312 then
	inst <= x"82242CB4";
end if;
if pc = 11316 then
	inst <= x"C43C0008";
end if;
if pc = 11320 then
	inst <= x"C17DFFFC";
end if;
if pc = 11324 then
	inst <= x"03DC0014";
end if;
if pc = 11328 then
	inst <= x"037E000C";
end if;
if pc = 11332 then
	inst <= x"C57DFFFC";
end if;
if pc = 11336 then
	inst <= x"82000794";
end if;
if pc = 11340 then
	inst <= x"07DC0014";
end if;
if pc = 11344 then
	inst <= x"0240FFFF";
end if;
if pc = 11348 then
	inst <= x"82242C88";
end if;
if pc = 11352 then
	inst <= x"02400003";
end if;
if pc = 11356 then
	inst <= x"C43C000C";
end if;
if pc = 11360 then
	inst <= x"C17DFFFC";
end if;
if pc = 11364 then
	inst <= x"00240000";
end if;
if pc = 11368 then
	inst <= x"03DC0018";
end if;
if pc = 11372 then
	inst <= x"037E000C";
end if;
if pc = 11376 then
	inst <= x"C57DFFFC";
end if;
if pc = 11380 then
	inst <= x"82002A44";
end if;
if pc = 11384 then
	inst <= x"07DC0018";
end if;
if pc = 11388 then
	inst <= x"C05C000C";
end if;
if pc = 11392 then
	inst <= x"C4420008";
end if;
if pc = 11396 then
	inst <= x"82002CA8";
end if;
if pc = 11400 then
	inst <= x"02200003";
end if;
if pc = 11404 then
	inst <= x"0240FFFF";
end if;
if pc = 11408 then
	inst <= x"C17DFFFC";
end if;
if pc = 11412 then
	inst <= x"03DC0018";
end if;
if pc = 11416 then
	inst <= x"037E000C";
end if;
if pc = 11420 then
	inst <= x"C57DFFFC";
end if;
if pc = 11424 then
	inst <= x"8200081C";
end if;
if pc = 11428 then
	inst <= x"07DC0018";
end if;
if pc = 11432 then
	inst <= x"C05C0008";
end if;
if pc = 11436 then
	inst <= x"C4420004";
end if;
if pc = 11440 then
	inst <= x"82002CD4";
end if;
if pc = 11444 then
	inst <= x"02200002";
end if;
if pc = 11448 then
	inst <= x"0240FFFF";
end if;
if pc = 11452 then
	inst <= x"C17DFFFC";
end if;
if pc = 11456 then
	inst <= x"03DC0018";
end if;
if pc = 11460 then
	inst <= x"037E000C";
end if;
if pc = 11464 then
	inst <= x"C57DFFFC";
end if;
if pc = 11468 then
	inst <= x"8200081C";
end if;
if pc = 11472 then
	inst <= x"07DC0018";
end if;
if pc = 11476 then
	inst <= x"C05C0004";
end if;
if pc = 11480 then
	inst <= x"C4420000";
end if;
if pc = 11484 then
	inst <= x"00420000";
end if;
if pc = 11488 then
	inst <= x"82002D08";
end if;
if pc = 11492 then
	inst <= x"02200001";
end if;
if pc = 11496 then
	inst <= x"0240FFFF";
end if;
if pc = 11500 then
	inst <= x"C17DFFFC";
end if;
if pc = 11504 then
	inst <= x"03DC0018";
end if;
if pc = 11508 then
	inst <= x"037E000C";
end if;
if pc = 11512 then
	inst <= x"C57DFFFC";
end if;
if pc = 11516 then
	inst <= x"8200081C";
end if;
if pc = 11520 then
	inst <= x"07DC0018";
end if;
if pc = 11524 then
	inst <= x"00420000";
end if;
if pc = 11528 then
	inst <= x"C0240000";
end if;
if pc = 11532 then
	inst <= x"0260FFFF";
end if;
if pc = 11536 then
	inst <= x"82262E68";
end if;
if pc = 11540 then
	inst <= x"C03C0000";
end if;
if pc = 11544 then
	inst <= x"02620001";
end if;
if pc = 11548 then
	inst <= x"C45C0010";
end if;
if pc = 11552 then
	inst <= x"C47C0014";
end if;
if pc = 11556 then
	inst <= x"C17DFFFC";
end if;
if pc = 11560 then
	inst <= x"03DC0020";
end if;
if pc = 11564 then
	inst <= x"037E000C";
end if;
if pc = 11568 then
	inst <= x"C57DFFFC";
end if;
if pc = 11572 then
	inst <= x"82000794";
end if;
if pc = 11576 then
	inst <= x"07DC0020";
end if;
if pc = 11580 then
	inst <= x"0240FFFF";
end if;
if pc = 11584 then
	inst <= x"82242DC8";
end if;
if pc = 11588 then
	inst <= x"C43C0018";
end if;
if pc = 11592 then
	inst <= x"C17DFFFC";
end if;
if pc = 11596 then
	inst <= x"03DC0024";
end if;
if pc = 11600 then
	inst <= x"037E000C";
end if;
if pc = 11604 then
	inst <= x"C57DFFFC";
end if;
if pc = 11608 then
	inst <= x"82000794";
end if;
if pc = 11612 then
	inst <= x"07DC0024";
end if;
if pc = 11616 then
	inst <= x"0240FFFF";
end if;
if pc = 11620 then
	inst <= x"82242D98";
end if;
if pc = 11624 then
	inst <= x"02400002";
end if;
if pc = 11628 then
	inst <= x"C43C001C";
end if;
if pc = 11632 then
	inst <= x"C17DFFFC";
end if;
if pc = 11636 then
	inst <= x"00240000";
end if;
if pc = 11640 then
	inst <= x"03DC0028";
end if;
if pc = 11644 then
	inst <= x"037E000C";
end if;
if pc = 11648 then
	inst <= x"C57DFFFC";
end if;
if pc = 11652 then
	inst <= x"82002A44";
end if;
if pc = 11656 then
	inst <= x"07DC0028";
end if;
if pc = 11660 then
	inst <= x"C05C001C";
end if;
if pc = 11664 then
	inst <= x"C4420004";
end if;
if pc = 11668 then
	inst <= x"82002DB8";
end if;
if pc = 11672 then
	inst <= x"02200002";
end if;
if pc = 11676 then
	inst <= x"0240FFFF";
end if;
if pc = 11680 then
	inst <= x"C17DFFFC";
end if;
if pc = 11684 then
	inst <= x"03DC0028";
end if;
if pc = 11688 then
	inst <= x"037E000C";
end if;
if pc = 11692 then
	inst <= x"C57DFFFC";
end if;
if pc = 11696 then
	inst <= x"8200081C";
end if;
if pc = 11700 then
	inst <= x"07DC0028";
end if;
if pc = 11704 then
	inst <= x"C05C0018";
end if;
if pc = 11708 then
	inst <= x"C4420000";
end if;
if pc = 11712 then
	inst <= x"00420000";
end if;
if pc = 11716 then
	inst <= x"82002DEC";
end if;
if pc = 11720 then
	inst <= x"02200001";
end if;
if pc = 11724 then
	inst <= x"0240FFFF";
end if;
if pc = 11728 then
	inst <= x"C17DFFFC";
end if;
if pc = 11732 then
	inst <= x"03DC0028";
end if;
if pc = 11736 then
	inst <= x"037E000C";
end if;
if pc = 11740 then
	inst <= x"C57DFFFC";
end if;
if pc = 11744 then
	inst <= x"8200081C";
end if;
if pc = 11748 then
	inst <= x"07DC0028";
end if;
if pc = 11752 then
	inst <= x"00420000";
end if;
if pc = 11756 then
	inst <= x"C0240000";
end if;
if pc = 11760 then
	inst <= x"0260FFFF";
end if;
if pc = 11764 then
	inst <= x"82262E34";
end if;
if pc = 11768 then
	inst <= x"C03C0014";
end if;
if pc = 11772 then
	inst <= x"02620001";
end if;
if pc = 11776 then
	inst <= x"C45C0020";
end if;
if pc = 11780 then
	inst <= x"C17DFFFC";
end if;
if pc = 11784 then
	inst <= x"00260000";
end if;
if pc = 11788 then
	inst <= x"03DC002C";
end if;
if pc = 11792 then
	inst <= x"037E000C";
end if;
if pc = 11796 then
	inst <= x"C57DFFFC";
end if;
if pc = 11800 then
	inst <= x"82002BEC";
end if;
if pc = 11804 then
	inst <= x"07DC002C";
end if;
if pc = 11808 then
	inst <= x"C05C0014";
end if;
if pc = 11812 then
	inst <= x"22440220";
end if;
if pc = 11816 then
	inst <= x"C07C0020";
end if;
if pc = 11820 then
	inst <= x"D4624000";
end if;
if pc = 11824 then
	inst <= x"82002E54";
end if;
if pc = 11828 then
	inst <= x"C03C0014";
end if;
if pc = 11832 then
	inst <= x"02220001";
end if;
if pc = 11836 then
	inst <= x"C17DFFFC";
end if;
if pc = 11840 then
	inst <= x"03DC002C";
end if;
if pc = 11844 then
	inst <= x"037E000C";
end if;
if pc = 11848 then
	inst <= x"C57DFFFC";
end if;
if pc = 11852 then
	inst <= x"8200081C";
end if;
if pc = 11856 then
	inst <= x"07DC002C";
end if;
if pc = 11860 then
	inst <= x"C05C0000";
end if;
if pc = 11864 then
	inst <= x"22440220";
end if;
if pc = 11868 then
	inst <= x"C07C0010";
end if;
if pc = 11872 then
	inst <= x"D4624000";
end if;
if pc = 11876 then
	inst <= x"C1FDFFFC";
end if;
if pc = 11880 then
	inst <= x"C03C0000";
end if;
if pc = 11884 then
	inst <= x"02220001";
end if;
if pc = 11888 then
	inst <= x"8200081C";
end if;
if pc = 11892 then
	inst <= x"C43C0000";
end if;
if pc = 11896 then
	inst <= x"C17DFFFC";
end if;
if pc = 11900 then
	inst <= x"03DC000C";
end if;
if pc = 11904 then
	inst <= x"037E000C";
end if;
if pc = 11908 then
	inst <= x"C57DFFFC";
end if;
if pc = 11912 then
	inst <= x"82000794";
end if;
if pc = 11916 then
	inst <= x"07DC000C";
end if;
if pc = 11920 then
	inst <= x"0240FFFF";
end if;
if pc = 11924 then
	inst <= x"82242F68";
end if;
if pc = 11928 then
	inst <= x"C43C0004";
end if;
if pc = 11932 then
	inst <= x"C17DFFFC";
end if;
if pc = 11936 then
	inst <= x"03DC0010";
end if;
if pc = 11940 then
	inst <= x"037E000C";
end if;
if pc = 11944 then
	inst <= x"C57DFFFC";
end if;
if pc = 11948 then
	inst <= x"82000794";
end if;
if pc = 11952 then
	inst <= x"07DC0010";
end if;
if pc = 11956 then
	inst <= x"0240FFFF";
end if;
if pc = 11960 then
	inst <= x"82242F3C";
end if;
if pc = 11964 then
	inst <= x"C43C0008";
end if;
if pc = 11968 then
	inst <= x"C17DFFFC";
end if;
if pc = 11972 then
	inst <= x"03DC0014";
end if;
if pc = 11976 then
	inst <= x"037E000C";
end if;
if pc = 11980 then
	inst <= x"C57DFFFC";
end if;
if pc = 11984 then
	inst <= x"82000794";
end if;
if pc = 11988 then
	inst <= x"07DC0014";
end if;
if pc = 11992 then
	inst <= x"0240FFFF";
end if;
if pc = 11996 then
	inst <= x"82242F10";
end if;
if pc = 12000 then
	inst <= x"02400003";
end if;
if pc = 12004 then
	inst <= x"C43C000C";
end if;
if pc = 12008 then
	inst <= x"C17DFFFC";
end if;
if pc = 12012 then
	inst <= x"00240000";
end if;
if pc = 12016 then
	inst <= x"03DC0018";
end if;
if pc = 12020 then
	inst <= x"037E000C";
end if;
if pc = 12024 then
	inst <= x"C57DFFFC";
end if;
if pc = 12028 then
	inst <= x"82002A44";
end if;
if pc = 12032 then
	inst <= x"07DC0018";
end if;
if pc = 12036 then
	inst <= x"C05C000C";
end if;
if pc = 12040 then
	inst <= x"C4420008";
end if;
if pc = 12044 then
	inst <= x"82002F30";
end if;
if pc = 12048 then
	inst <= x"02200003";
end if;
if pc = 12052 then
	inst <= x"0240FFFF";
end if;
if pc = 12056 then
	inst <= x"C17DFFFC";
end if;
if pc = 12060 then
	inst <= x"03DC0018";
end if;
if pc = 12064 then
	inst <= x"037E000C";
end if;
if pc = 12068 then
	inst <= x"C57DFFFC";
end if;
if pc = 12072 then
	inst <= x"8200081C";
end if;
if pc = 12076 then
	inst <= x"07DC0018";
end if;
if pc = 12080 then
	inst <= x"C05C0008";
end if;
if pc = 12084 then
	inst <= x"C4420004";
end if;
if pc = 12088 then
	inst <= x"82002F5C";
end if;
if pc = 12092 then
	inst <= x"02200002";
end if;
if pc = 12096 then
	inst <= x"0240FFFF";
end if;
if pc = 12100 then
	inst <= x"C17DFFFC";
end if;
if pc = 12104 then
	inst <= x"03DC0018";
end if;
if pc = 12108 then
	inst <= x"037E000C";
end if;
if pc = 12112 then
	inst <= x"C57DFFFC";
end if;
if pc = 12116 then
	inst <= x"8200081C";
end if;
if pc = 12120 then
	inst <= x"07DC0018";
end if;
if pc = 12124 then
	inst <= x"C05C0004";
end if;
if pc = 12128 then
	inst <= x"C4420000";
end if;
if pc = 12132 then
	inst <= x"82002F88";
end if;
if pc = 12136 then
	inst <= x"02200001";
end if;
if pc = 12140 then
	inst <= x"0240FFFF";
end if;
if pc = 12144 then
	inst <= x"C17DFFFC";
end if;
if pc = 12148 then
	inst <= x"03DC0018";
end if;
if pc = 12152 then
	inst <= x"037E000C";
end if;
if pc = 12156 then
	inst <= x"C57DFFFC";
end if;
if pc = 12160 then
	inst <= x"8200081C";
end if;
if pc = 12164 then
	inst <= x"07DC0018";
end if;
if pc = 12168 then
	inst <= x"C0420000";
end if;
if pc = 12172 then
	inst <= x"0260FFFF";
end if;
if pc = 12176 then
	inst <= x"82463178";
end if;
if pc = 12180 then
	inst <= x"024001E0";
end if;
if pc = 12184 then
	inst <= x"C07C0000";
end if;
if pc = 12188 then
	inst <= x"22860220";
end if;
if pc = 12192 then
	inst <= x"D4248000";
end if;
if pc = 12196 then
	inst <= x"02260001";
end if;
if pc = 12200 then
	inst <= x"C45C0010";
end if;
if pc = 12204 then
	inst <= x"C43C0014";
end if;
if pc = 12208 then
	inst <= x"C17DFFFC";
end if;
if pc = 12212 then
	inst <= x"03DC0020";
end if;
if pc = 12216 then
	inst <= x"037E000C";
end if;
if pc = 12220 then
	inst <= x"C57DFFFC";
end if;
if pc = 12224 then
	inst <= x"82000794";
end if;
if pc = 12228 then
	inst <= x"07DC0020";
end if;
if pc = 12232 then
	inst <= x"0240FFFF";
end if;
if pc = 12236 then
	inst <= x"82243050";
end if;
if pc = 12240 then
	inst <= x"C43C0018";
end if;
if pc = 12244 then
	inst <= x"C17DFFFC";
end if;
if pc = 12248 then
	inst <= x"03DC0024";
end if;
if pc = 12252 then
	inst <= x"037E000C";
end if;
if pc = 12256 then
	inst <= x"C57DFFFC";
end if;
if pc = 12260 then
	inst <= x"82000794";
end if;
if pc = 12264 then
	inst <= x"07DC0024";
end if;
if pc = 12268 then
	inst <= x"0240FFFF";
end if;
if pc = 12272 then
	inst <= x"82243024";
end if;
if pc = 12276 then
	inst <= x"02400002";
end if;
if pc = 12280 then
	inst <= x"C43C001C";
end if;
if pc = 12284 then
	inst <= x"C17DFFFC";
end if;
if pc = 12288 then
	inst <= x"00240000";
end if;
if pc = 12292 then
	inst <= x"03DC0028";
end if;
if pc = 12296 then
	inst <= x"037E000C";
end if;
if pc = 12300 then
	inst <= x"C57DFFFC";
end if;
if pc = 12304 then
	inst <= x"82002A44";
end if;
if pc = 12308 then
	inst <= x"07DC0028";
end if;
if pc = 12312 then
	inst <= x"C05C001C";
end if;
if pc = 12316 then
	inst <= x"C4420004";
end if;
if pc = 12320 then
	inst <= x"82003044";
end if;
if pc = 12324 then
	inst <= x"02200002";
end if;
if pc = 12328 then
	inst <= x"0240FFFF";
end if;
if pc = 12332 then
	inst <= x"C17DFFFC";
end if;
if pc = 12336 then
	inst <= x"03DC0028";
end if;
if pc = 12340 then
	inst <= x"037E000C";
end if;
if pc = 12344 then
	inst <= x"C57DFFFC";
end if;
if pc = 12348 then
	inst <= x"8200081C";
end if;
if pc = 12352 then
	inst <= x"07DC0028";
end if;
if pc = 12356 then
	inst <= x"C05C0018";
end if;
if pc = 12360 then
	inst <= x"C4420000";
end if;
if pc = 12364 then
	inst <= x"82003070";
end if;
if pc = 12368 then
	inst <= x"02200001";
end if;
if pc = 12372 then
	inst <= x"0240FFFF";
end if;
if pc = 12376 then
	inst <= x"C17DFFFC";
end if;
if pc = 12380 then
	inst <= x"03DC0028";
end if;
if pc = 12384 then
	inst <= x"037E000C";
end if;
if pc = 12388 then
	inst <= x"C57DFFFC";
end if;
if pc = 12392 then
	inst <= x"8200081C";
end if;
if pc = 12396 then
	inst <= x"07DC0028";
end if;
if pc = 12400 then
	inst <= x"C0420000";
end if;
if pc = 12404 then
	inst <= x"0260FFFF";
end if;
if pc = 12408 then
	inst <= x"82463174";
end if;
if pc = 12412 then
	inst <= x"C05C0014";
end if;
if pc = 12416 then
	inst <= x"22640220";
end if;
if pc = 12420 then
	inst <= x"C09C0010";
end if;
if pc = 12424 then
	inst <= x"D4286000";
end if;
if pc = 12428 then
	inst <= x"02240001";
end if;
if pc = 12432 then
	inst <= x"C43C0020";
end if;
if pc = 12436 then
	inst <= x"C17DFFFC";
end if;
if pc = 12440 then
	inst <= x"03DC002C";
end if;
if pc = 12444 then
	inst <= x"037E000C";
end if;
if pc = 12448 then
	inst <= x"C57DFFFC";
end if;
if pc = 12452 then
	inst <= x"82000794";
end if;
if pc = 12456 then
	inst <= x"07DC002C";
end if;
if pc = 12460 then
	inst <= x"0240FFFF";
end if;
if pc = 12464 then
	inst <= x"822430E4";
end if;
if pc = 12468 then
	inst <= x"02400001";
end if;
if pc = 12472 then
	inst <= x"C43C0024";
end if;
if pc = 12476 then
	inst <= x"C17DFFFC";
end if;
if pc = 12480 then
	inst <= x"00240000";
end if;
if pc = 12484 then
	inst <= x"03DC0030";
end if;
if pc = 12488 then
	inst <= x"037E000C";
end if;
if pc = 12492 then
	inst <= x"C57DFFFC";
end if;
if pc = 12496 then
	inst <= x"82002A44";
end if;
if pc = 12500 then
	inst <= x"07DC0030";
end if;
if pc = 12504 then
	inst <= x"C05C0024";
end if;
if pc = 12508 then
	inst <= x"C4420000";
end if;
if pc = 12512 then
	inst <= x"82003104";
end if;
if pc = 12516 then
	inst <= x"02200001";
end if;
if pc = 12520 then
	inst <= x"0240FFFF";
end if;
if pc = 12524 then
	inst <= x"C17DFFFC";
end if;
if pc = 12528 then
	inst <= x"03DC0030";
end if;
if pc = 12532 then
	inst <= x"037E000C";
end if;
if pc = 12536 then
	inst <= x"C57DFFFC";
end if;
if pc = 12540 then
	inst <= x"8200081C";
end if;
if pc = 12544 then
	inst <= x"07DC0030";
end if;
if pc = 12548 then
	inst <= x"C0420000";
end if;
if pc = 12552 then
	inst <= x"0260FFFF";
end if;
if pc = 12556 then
	inst <= x"82463170";
end if;
if pc = 12560 then
	inst <= x"C05C0020";
end if;
if pc = 12564 then
	inst <= x"22640220";
end if;
if pc = 12568 then
	inst <= x"C09C0010";
end if;
if pc = 12572 then
	inst <= x"D4286000";
end if;
if pc = 12576 then
	inst <= x"02240001";
end if;
if pc = 12580 then
	inst <= x"02400000";
end if;
if pc = 12584 then
	inst <= x"C43C0028";
end if;
if pc = 12588 then
	inst <= x"C17DFFFC";
end if;
if pc = 12592 then
	inst <= x"00240000";
end if;
if pc = 12596 then
	inst <= x"03DC0034";
end if;
if pc = 12600 then
	inst <= x"037E000C";
end if;
if pc = 12604 then
	inst <= x"C57DFFFC";
end if;
if pc = 12608 then
	inst <= x"82002A44";
end if;
if pc = 12612 then
	inst <= x"07DC0034";
end if;
if pc = 12616 then
	inst <= x"C0420000";
end if;
if pc = 12620 then
	inst <= x"0260FFFF";
end if;
if pc = 12624 then
	inst <= x"8246316C";
end if;
if pc = 12628 then
	inst <= x"C05C0028";
end if;
if pc = 12632 then
	inst <= x"22640220";
end if;
if pc = 12636 then
	inst <= x"C09C0010";
end if;
if pc = 12640 then
	inst <= x"D4286000";
end if;
if pc = 12644 then
	inst <= x"02240001";
end if;
if pc = 12648 then
	inst <= x"82002E74";
end if;
if pc = 12652 then
	inst <= x"C1FDFFFC";
end if;
if pc = 12656 then
	inst <= x"C1FDFFFC";
end if;
if pc = 12660 then
	inst <= x"C1FDFFFC";
end if;
if pc = 12664 then
	inst <= x"C1FDFFFC";
end if;
if pc = 12668 then
	inst <= x"22C60220";
end if;
if pc = 12672 then
	inst <= x"D884C000";
end if;
if pc = 12676 then
	inst <= x"8A80329C";
end if;
if pc = 12680 then
	inst <= x"C0C20010";
end if;
if pc = 12684 then
	inst <= x"C0220018";
end if;
if pc = 12688 then
	inst <= x"8E80319C";
end if;
if pc = 12692 then
	inst <= x"02E00000";
end if;
if pc = 12696 then
	inst <= x"820031A0";
end if;
if pc = 12700 then
	inst <= x"02E00001";
end if;
if pc = 12704 then
	inst <= x"822031B8";
end if;
if pc = 12708 then
	inst <= x"8E8031B0";
end if;
if pc = 12712 then
	inst <= x"02200001";
end if;
if pc = 12716 then
	inst <= x"820031B4";
end if;
if pc = 12720 then
	inst <= x"02200000";
end if;
if pc = 12724 then
	inst <= x"820031BC";
end if;
if pc = 12728 then
	inst <= x"002E0000";
end if;
if pc = 12732 then
	inst <= x"22660220";
end if;
if pc = 12736 then
	inst <= x"D8AC6000";
end if;
if pc = 12740 then
	inst <= x"822031CC";
end if;
if pc = 12744 then
	inst <= x"820031D0";
end if;
if pc = 12748 then
	inst <= x"44A0A000";
end if;
if pc = 12752 then
	inst <= x"442A2000";
end if;
if pc = 12756 then
	inst <= x"CC7C0000";
end if;
if pc = 12760 then
	inst <= x"C4BC0008";
end if;
if pc = 12764 then
	inst <= x"C4DC000C";
end if;
if pc = 12768 then
	inst <= x"CC5C0010";
end if;
if pc = 12772 then
	inst <= x"C45C0018";
end if;
if pc = 12776 then
	inst <= x"C49C001C";
end if;
if pc = 12780 then
	inst <= x"CC3C0020";
end if;
if pc = 12784 then
	inst <= x"C17DFFFC";
end if;
if pc = 12788 then
	inst <= x"40208000";
end if;
if pc = 12792 then
	inst <= x"03DC0030";
end if;
if pc = 12796 then
	inst <= x"037E000C";
end if;
if pc = 12800 then
	inst <= x"C57DFFFC";
end if;
if pc = 12804 then
	inst <= x"82000844";
end if;
if pc = 12808 then
	inst <= x"07DC0030";
end if;
if pc = 12812 then
	inst <= x"C85C0020";
end if;
if pc = 12816 then
	inst <= x"48242000";
end if;
if pc = 12820 then
	inst <= x"C03C001C";
end if;
if pc = 12824 then
	inst <= x"22420220";
end if;
if pc = 12828 then
	inst <= x"C07C0018";
end if;
if pc = 12832 then
	inst <= x"D8464000";
end if;
if pc = 12836 then
	inst <= x"48424000";
end if;
if pc = 12840 then
	inst <= x"C87C0010";
end if;
if pc = 12844 then
	inst <= x"40446000";
end if;
if pc = 12848 then
	inst <= x"8E403238";
end if;
if pc = 12852 then
	inst <= x"8200323C";
end if;
if pc = 12856 then
	inst <= x"44404000";
end if;
if pc = 12860 then
	inst <= x"22220220";
end if;
if pc = 12864 then
	inst <= x"C05C000C";
end if;
if pc = 12868 then
	inst <= x"D8642000";
end if;
if pc = 12872 then
	inst <= x"8E463254";
end if;
if pc = 12876 then
	inst <= x"02200000";
end if;
if pc = 12880 then
	inst <= x"C1FDFFFC";
end if;
if pc = 12884 then
	inst <= x"C03C0008";
end if;
if pc = 12888 then
	inst <= x"22820220";
end if;
if pc = 12892 then
	inst <= x"D8468000";
end if;
if pc = 12896 then
	inst <= x"48424000";
end if;
if pc = 12900 then
	inst <= x"C87C0000";
end if;
if pc = 12904 then
	inst <= x"40446000";
end if;
if pc = 12908 then
	inst <= x"8E403274";
end if;
if pc = 12912 then
	inst <= x"82003278";
end if;
if pc = 12916 then
	inst <= x"44404000";
end if;
if pc = 12920 then
	inst <= x"22220220";
end if;
if pc = 12924 then
	inst <= x"D8642000";
end if;
if pc = 12928 then
	inst <= x"8E46328C";
end if;
if pc = 12932 then
	inst <= x"02200000";
end if;
if pc = 12936 then
	inst <= x"C1FDFFFC";
end if;
if pc = 12940 then
	inst <= x"022002AC";
end if;
if pc = 12944 then
	inst <= x"CC220000";
end if;
if pc = 12948 then
	inst <= x"02200001";
end if;
if pc = 12952 then
	inst <= x"C1FDFFFC";
end if;
if pc = 12956 then
	inst <= x"02200000";
end if;
if pc = 12960 then
	inst <= x"C1FDFFFC";
end if;
if pc = 12964 then
	inst <= x"C0220010";
end if;
if pc = 12968 then
	inst <= x"C8840000";
end if;
if pc = 12972 then
	inst <= x"C8A20000";
end if;
if pc = 12976 then
	inst <= x"4888A000";
end if;
if pc = 12980 then
	inst <= x"C8A40004";
end if;
if pc = 12984 then
	inst <= x"C8C20004";
end if;
if pc = 12988 then
	inst <= x"48AAC000";
end if;
if pc = 12992 then
	inst <= x"4088A000";
end if;
if pc = 12996 then
	inst <= x"C8A40008";
end if;
if pc = 13000 then
	inst <= x"C8C20008";
end if;
if pc = 13004 then
	inst <= x"48AAC000";
end if;
if pc = 13008 then
	inst <= x"4088A000";
end if;
if pc = 13012 then
	inst <= x"8E0832E0";
end if;
if pc = 13016 then
	inst <= x"02200000";
end if;
if pc = 13020 then
	inst <= x"C1FDFFFC";
end if;
if pc = 13024 then
	inst <= x"024002AC";
end if;
if pc = 13028 then
	inst <= x"C8A20000";
end if;
if pc = 13032 then
	inst <= x"482A2000";
end if;
if pc = 13036 then
	inst <= x"C8A20004";
end if;
if pc = 13040 then
	inst <= x"484A4000";
end if;
if pc = 13044 then
	inst <= x"40224000";
end if;
if pc = 13048 then
	inst <= x"C8420008";
end if;
if pc = 13052 then
	inst <= x"48446000";
end if;
if pc = 13056 then
	inst <= x"40224000";
end if;
if pc = 13060 then
	inst <= x"44202000";
end if;
if pc = 13064 then
	inst <= x"C45C0000";
end if;
if pc = 13068 then
	inst <= x"CC3C0008";
end if;
if pc = 13072 then
	inst <= x"C17DFFFC";
end if;
if pc = 13076 then
	inst <= x"40208000";
end if;
if pc = 13080 then
	inst <= x"03DC0018";
end if;
if pc = 13084 then
	inst <= x"037E000C";
end if;
if pc = 13088 then
	inst <= x"C57DFFFC";
end if;
if pc = 13092 then
	inst <= x"82000844";
end if;
if pc = 13096 then
	inst <= x"07DC0018";
end if;
if pc = 13100 then
	inst <= x"C85C0008";
end if;
if pc = 13104 then
	inst <= x"48242000";
end if;
if pc = 13108 then
	inst <= x"C03C0000";
end if;
if pc = 13112 then
	inst <= x"CC220000";
end if;
if pc = 13116 then
	inst <= x"02200001";
end if;
if pc = 13120 then
	inst <= x"C1FDFFFC";
end if;
if pc = 13124 then
	inst <= x"48822000";
end if;
if pc = 13128 then
	inst <= x"C0420010";
end if;
if pc = 13132 then
	inst <= x"C8A40000";
end if;
if pc = 13136 then
	inst <= x"4888A000";
end if;
if pc = 13140 then
	inst <= x"48A44000";
end if;
if pc = 13144 then
	inst <= x"C0420010";
end if;
if pc = 13148 then
	inst <= x"C8C40004";
end if;
if pc = 13152 then
	inst <= x"48AAC000";
end if;
if pc = 13156 then
	inst <= x"4088A000";
end if;
if pc = 13160 then
	inst <= x"48A66000";
end if;
if pc = 13164 then
	inst <= x"C0420010";
end if;
if pc = 13168 then
	inst <= x"C8C40008";
end if;
if pc = 13172 then
	inst <= x"48AAC000";
end if;
if pc = 13176 then
	inst <= x"4088A000";
end if;
if pc = 13180 then
	inst <= x"C042000C";
end if;
if pc = 13184 then
	inst <= x"824033C4";
end if;
if pc = 13188 then
	inst <= x"48A46000";
end if;
if pc = 13192 then
	inst <= x"C0420024";
end if;
if pc = 13196 then
	inst <= x"C8C40000";
end if;
if pc = 13200 then
	inst <= x"48AAC000";
end if;
if pc = 13204 then
	inst <= x"4088A000";
end if;
if pc = 13208 then
	inst <= x"48662000";
end if;
if pc = 13212 then
	inst <= x"C0420024";
end if;
if pc = 13216 then
	inst <= x"C8A40004";
end if;
if pc = 13220 then
	inst <= x"4866A000";
end if;
if pc = 13224 then
	inst <= x"40686000";
end if;
if pc = 13228 then
	inst <= x"48224000";
end if;
if pc = 13232 then
	inst <= x"C0220024";
end if;
if pc = 13236 then
	inst <= x"C8420008";
end if;
if pc = 13240 then
	inst <= x"48224000";
end if;
if pc = 13244 then
	inst <= x"40262000";
end if;
if pc = 13248 then
	inst <= x"C1FDFFFC";
end if;
if pc = 13252 then
	inst <= x"40208000";
end if;
if pc = 13256 then
	inst <= x"C1FDFFFC";
end if;
if pc = 13260 then
	inst <= x"48E28000";
end if;
if pc = 13264 then
	inst <= x"C0420010";
end if;
if pc = 13268 then
	inst <= x"C9040000";
end if;
if pc = 13272 then
	inst <= x"48EF0000";
end if;
if pc = 13276 then
	inst <= x"4904A000";
end if;
if pc = 13280 then
	inst <= x"C0420010";
end if;
if pc = 13284 then
	inst <= x"C9240004";
end if;
if pc = 13288 then
	inst <= x"49112000";
end if;
if pc = 13292 then
	inst <= x"40EF0000";
end if;
if pc = 13296 then
	inst <= x"4906C000";
end if;
if pc = 13300 then
	inst <= x"C0420010";
end if;
if pc = 13304 then
	inst <= x"C9240008";
end if;
if pc = 13308 then
	inst <= x"49112000";
end if;
if pc = 13312 then
	inst <= x"40EF0000";
end if;
if pc = 13316 then
	inst <= x"C042000C";
end if;
if pc = 13320 then
	inst <= x"82403498";
end if;
if pc = 13324 then
	inst <= x"4906A000";
end if;
if pc = 13328 then
	inst <= x"4924C000";
end if;
if pc = 13332 then
	inst <= x"41112000";
end if;
if pc = 13336 then
	inst <= x"C0420024";
end if;
if pc = 13340 then
	inst <= x"C9240000";
end if;
if pc = 13344 then
	inst <= x"49112000";
end if;
if pc = 13348 then
	inst <= x"48C2C000";
end if;
if pc = 13352 then
	inst <= x"48668000";
end if;
if pc = 13356 then
	inst <= x"406C6000";
end if;
if pc = 13360 then
	inst <= x"C0420024";
end if;
if pc = 13364 then
	inst <= x"C8C40004";
end if;
if pc = 13368 then
	inst <= x"4866C000";
end if;
if pc = 13372 then
	inst <= x"40706000";
end if;
if pc = 13376 then
	inst <= x"4822A000";
end if;
if pc = 13380 then
	inst <= x"48448000";
end if;
if pc = 13384 then
	inst <= x"40224000";
end if;
if pc = 13388 then
	inst <= x"C0220024";
end if;
if pc = 13392 then
	inst <= x"C8420008";
end if;
if pc = 13396 then
	inst <= x"48224000";
end if;
if pc = 13400 then
	inst <= x"40262000";
end if;
if pc = 13404 then
	inst <= x"C8400080";
end if;
if pc = 13408 then
	inst <= x"CCFC0000";
end if;
if pc = 13412 then
	inst <= x"CC3C0008";
end if;
if pc = 13416 then
	inst <= x"C17DFFFC";
end if;
if pc = 13420 then
	inst <= x"40204000";
end if;
if pc = 13424 then
	inst <= x"03DC0018";
end if;
if pc = 13428 then
	inst <= x"037E000C";
end if;
if pc = 13432 then
	inst <= x"C57DFFFC";
end if;
if pc = 13436 then
	inst <= x"82000844";
end if;
if pc = 13440 then
	inst <= x"07DC0018";
end if;
if pc = 13444 then
	inst <= x"C85C0008";
end if;
if pc = 13448 then
	inst <= x"48242000";
end if;
if pc = 13452 then
	inst <= x"C85C0000";
end if;
if pc = 13456 then
	inst <= x"40242000";
end if;
if pc = 13460 then
	inst <= x"C1FDFFFC";
end if;
if pc = 13464 then
	inst <= x"4020E000";
end if;
if pc = 13468 then
	inst <= x"C1FDFFFC";
end if;
if pc = 13472 then
	inst <= x"C8840000";
end if;
if pc = 13476 then
	inst <= x"C8A40004";
end if;
if pc = 13480 then
	inst <= x"C8C40008";
end if;
if pc = 13484 then
	inst <= x"48E88000";
end if;
if pc = 13488 then
	inst <= x"C0620010";
end if;
if pc = 13492 then
	inst <= x"C9060000";
end if;
if pc = 13496 then
	inst <= x"48EF0000";
end if;
if pc = 13500 then
	inst <= x"490AA000";
end if;
if pc = 13504 then
	inst <= x"C0620010";
end if;
if pc = 13508 then
	inst <= x"C9260004";
end if;
if pc = 13512 then
	inst <= x"49112000";
end if;
if pc = 13516 then
	inst <= x"40EF0000";
end if;
if pc = 13520 then
	inst <= x"490CC000";
end if;
if pc = 13524 then
	inst <= x"C0620010";
end if;
if pc = 13528 then
	inst <= x"C9260008";
end if;
if pc = 13532 then
	inst <= x"49112000";
end if;
if pc = 13536 then
	inst <= x"40EF0000";
end if;
if pc = 13540 then
	inst <= x"C062000C";
end if;
if pc = 13544 then
	inst <= x"8260352C";
end if;
if pc = 13548 then
	inst <= x"490AC000";
end if;
if pc = 13552 then
	inst <= x"C0620024";
end if;
if pc = 13556 then
	inst <= x"C9260000";
end if;
if pc = 13560 then
	inst <= x"49112000";
end if;
if pc = 13564 then
	inst <= x"40EF0000";
end if;
if pc = 13568 then
	inst <= x"48CC8000";
end if;
if pc = 13572 then
	inst <= x"C0620024";
end if;
if pc = 13576 then
	inst <= x"C9060004";
end if;
if pc = 13580 then
	inst <= x"48CD0000";
end if;
if pc = 13584 then
	inst <= x"40CEC000";
end if;
if pc = 13588 then
	inst <= x"4888A000";
end if;
if pc = 13592 then
	inst <= x"C0620024";
end if;
if pc = 13596 then
	inst <= x"C8A60008";
end if;
if pc = 13600 then
	inst <= x"4888A000";
end if;
if pc = 13604 then
	inst <= x"408C8000";
end if;
if pc = 13608 then
	inst <= x"82003530";
end if;
if pc = 13612 then
	inst <= x"4080E000";
end if;
if pc = 13616 then
	inst <= x"8A8036CC";
end if;
if pc = 13620 then
	inst <= x"C8A40000";
end if;
if pc = 13624 then
	inst <= x"C8C40004";
end if;
if pc = 13628 then
	inst <= x"C8E40008";
end if;
if pc = 13632 then
	inst <= x"CC9C0000";
end if;
if pc = 13636 then
	inst <= x"CC7C0008";
end if;
if pc = 13640 then
	inst <= x"CC5C0010";
end if;
if pc = 13644 then
	inst <= x"C43C0018";
end if;
if pc = 13648 then
	inst <= x"CC3C0020";
end if;
if pc = 13652 then
	inst <= x"C17DFFFC";
end if;
if pc = 13656 then
	inst <= x"40802000";
end if;
if pc = 13660 then
	inst <= x"4020A000";
end if;
if pc = 13664 then
	inst <= x"40A04000";
end if;
if pc = 13668 then
	inst <= x"4040C000";
end if;
if pc = 13672 then
	inst <= x"40C06000";
end if;
if pc = 13676 then
	inst <= x"4060E000";
end if;
if pc = 13680 then
	inst <= x"03DC0030";
end if;
if pc = 13684 then
	inst <= x"037E000C";
end if;
if pc = 13688 then
	inst <= x"C57DFFFC";
end if;
if pc = 13692 then
	inst <= x"820033CC";
end if;
if pc = 13696 then
	inst <= x"07DC0030";
end if;
if pc = 13700 then
	inst <= x"C85C0020";
end if;
if pc = 13704 then
	inst <= x"48644000";
end if;
if pc = 13708 then
	inst <= x"C03C0018";
end if;
if pc = 13712 then
	inst <= x"C0420010";
end if;
if pc = 13716 then
	inst <= x"C8840000";
end if;
if pc = 13720 then
	inst <= x"48668000";
end if;
if pc = 13724 then
	inst <= x"C89C0010";
end if;
if pc = 13728 then
	inst <= x"48A88000";
end if;
if pc = 13732 then
	inst <= x"C0420010";
end if;
if pc = 13736 then
	inst <= x"C8C40004";
end if;
if pc = 13740 then
	inst <= x"48AAC000";
end if;
if pc = 13744 then
	inst <= x"4066A000";
end if;
if pc = 13748 then
	inst <= x"C8BC0008";
end if;
if pc = 13752 then
	inst <= x"48CAA000";
end if;
if pc = 13756 then
	inst <= x"C0420010";
end if;
if pc = 13760 then
	inst <= x"C8E40008";
end if;
if pc = 13764 then
	inst <= x"48CCE000";
end if;
if pc = 13768 then
	inst <= x"4066C000";
end if;
if pc = 13772 then
	inst <= x"C042000C";
end if;
if pc = 13776 then
	inst <= x"82403614";
end if;
if pc = 13780 then
	inst <= x"48C8A000";
end if;
if pc = 13784 then
	inst <= x"C0420024";
end if;
if pc = 13788 then
	inst <= x"C8E40000";
end if;
if pc = 13792 then
	inst <= x"48CCE000";
end if;
if pc = 13796 then
	inst <= x"4066C000";
end if;
if pc = 13800 then
	inst <= x"48AA4000";
end if;
if pc = 13804 then
	inst <= x"C0420024";
end if;
if pc = 13808 then
	inst <= x"C8C40004";
end if;
if pc = 13812 then
	inst <= x"48AAC000";
end if;
if pc = 13816 then
	inst <= x"4066A000";
end if;
if pc = 13820 then
	inst <= x"48448000";
end if;
if pc = 13824 then
	inst <= x"C0420024";
end if;
if pc = 13828 then
	inst <= x"C8840008";
end if;
if pc = 13832 then
	inst <= x"48448000";
end if;
if pc = 13836 then
	inst <= x"40464000";
end if;
if pc = 13840 then
	inst <= x"82003618";
end if;
if pc = 13844 then
	inst <= x"40406000";
end if;
if pc = 13848 then
	inst <= x"C0420004";
end if;
if pc = 13852 then
	inst <= x"02600003";
end if;
if pc = 13856 then
	inst <= x"82463628";
end if;
if pc = 13860 then
	inst <= x"82003630";
end if;
if pc = 13864 then
	inst <= x"C86000A8";
end if;
if pc = 13868 then
	inst <= x"44446000";
end if;
if pc = 13872 then
	inst <= x"48622000";
end if;
if pc = 13876 then
	inst <= x"C89C0000";
end if;
if pc = 13880 then
	inst <= x"48484000";
end if;
if pc = 13884 then
	inst <= x"44464000";
end if;
if pc = 13888 then
	inst <= x"8E04364C";
end if;
if pc = 13892 then
	inst <= x"02200000";
end if;
if pc = 13896 then
	inst <= x"C1FDFFFC";
end if;
if pc = 13900 then
	inst <= x"CC3C0028";
end if;
if pc = 13904 then
	inst <= x"C17DFFFC";
end if;
if pc = 13908 then
	inst <= x"40204000";
end if;
if pc = 13912 then
	inst <= x"03DC0038";
end if;
if pc = 13916 then
	inst <= x"037E000C";
end if;
if pc = 13920 then
	inst <= x"C57DFFFC";
end if;
if pc = 13924 then
	inst <= x"8200083C";
end if;
if pc = 13928 then
	inst <= x"07DC0038";
end if;
if pc = 13932 then
	inst <= x"C03C0018";
end if;
if pc = 13936 then
	inst <= x"C0220018";
end if;
if pc = 13940 then
	inst <= x"8220367C";
end if;
if pc = 13944 then
	inst <= x"82003680";
end if;
if pc = 13948 then
	inst <= x"44202000";
end if;
if pc = 13952 then
	inst <= x"022002AC";
end if;
if pc = 13956 then
	inst <= x"C85C0028";
end if;
if pc = 13960 then
	inst <= x"44224000";
end if;
if pc = 13964 then
	inst <= x"C85C0000";
end if;
if pc = 13968 then
	inst <= x"C43C0030";
end if;
if pc = 13972 then
	inst <= x"CC3C0038";
end if;
if pc = 13976 then
	inst <= x"C17DFFFC";
end if;
if pc = 13980 then
	inst <= x"40204000";
end if;
if pc = 13984 then
	inst <= x"03DC0048";
end if;
if pc = 13988 then
	inst <= x"037E000C";
end if;
if pc = 13992 then
	inst <= x"C57DFFFC";
end if;
if pc = 13996 then
	inst <= x"82000844";
end if;
if pc = 14000 then
	inst <= x"07DC0048";
end if;
if pc = 14004 then
	inst <= x"C85C0038";
end if;
if pc = 14008 then
	inst <= x"48242000";
end if;
if pc = 14012 then
	inst <= x"C03C0030";
end if;
if pc = 14016 then
	inst <= x"CC220000";
end if;
if pc = 14020 then
	inst <= x"02200001";
end if;
if pc = 14024 then
	inst <= x"C1FDFFFC";
end if;
if pc = 14028 then
	inst <= x"02200000";
end if;
if pc = 14032 then
	inst <= x"C1FDFFFC";
end if;
if pc = 14036 then
	inst <= x"028000C8";
end if;
if pc = 14040 then
	inst <= x"22220220";
end if;
if pc = 14044 then
	inst <= x"D0282000";
end if;
if pc = 14048 then
	inst <= x"C8260000";
end if;
if pc = 14052 then
	inst <= x"C0820014";
end if;
if pc = 14056 then
	inst <= x"C8480000";
end if;
if pc = 14060 then
	inst <= x"44224000";
end if;
if pc = 14064 then
	inst <= x"C8460004";
end if;
if pc = 14068 then
	inst <= x"C0820014";
end if;
if pc = 14072 then
	inst <= x"C8680004";
end if;
if pc = 14076 then
	inst <= x"44446000";
end if;
if pc = 14080 then
	inst <= x"C8660008";
end if;
if pc = 14084 then
	inst <= x"C0620014";
end if;
if pc = 14088 then
	inst <= x"C8860008";
end if;
if pc = 14092 then
	inst <= x"44668000";
end if;
if pc = 14096 then
	inst <= x"C0620004";
end if;
if pc = 14100 then
	inst <= x"02800001";
end if;
if pc = 14104 then
	inst <= x"826837C8";
end if;
if pc = 14108 then
	inst <= x"02800002";
end if;
if pc = 14112 then
	inst <= x"82683728";
end if;
if pc = 14116 then
	inst <= x"820034A0";
end if;
if pc = 14120 then
	inst <= x"C0220010";
end if;
if pc = 14124 then
	inst <= x"C8840000";
end if;
if pc = 14128 then
	inst <= x"C8A20000";
end if;
if pc = 14132 then
	inst <= x"4888A000";
end if;
if pc = 14136 then
	inst <= x"C8A40004";
end if;
if pc = 14140 then
	inst <= x"C8C20004";
end if;
if pc = 14144 then
	inst <= x"48AAC000";
end if;
if pc = 14148 then
	inst <= x"4088A000";
end if;
if pc = 14152 then
	inst <= x"C8A40008";
end if;
if pc = 14156 then
	inst <= x"C8C20008";
end if;
if pc = 14160 then
	inst <= x"48AAC000";
end if;
if pc = 14164 then
	inst <= x"4088A000";
end if;
if pc = 14168 then
	inst <= x"8E083764";
end if;
if pc = 14172 then
	inst <= x"02200000";
end if;
if pc = 14176 then
	inst <= x"C1FDFFFC";
end if;
if pc = 14180 then
	inst <= x"024002AC";
end if;
if pc = 14184 then
	inst <= x"C8A20000";
end if;
if pc = 14188 then
	inst <= x"482A2000";
end if;
if pc = 14192 then
	inst <= x"C8A20004";
end if;
if pc = 14196 then
	inst <= x"484A4000";
end if;
if pc = 14200 then
	inst <= x"40224000";
end if;
if pc = 14204 then
	inst <= x"C8420008";
end if;
if pc = 14208 then
	inst <= x"48446000";
end if;
if pc = 14212 then
	inst <= x"40224000";
end if;
if pc = 14216 then
	inst <= x"44202000";
end if;
if pc = 14220 then
	inst <= x"C45C0000";
end if;
if pc = 14224 then
	inst <= x"CC3C0008";
end if;
if pc = 14228 then
	inst <= x"C17DFFFC";
end if;
if pc = 14232 then
	inst <= x"40208000";
end if;
if pc = 14236 then
	inst <= x"03DC0018";
end if;
if pc = 14240 then
	inst <= x"037E000C";
end if;
if pc = 14244 then
	inst <= x"C57DFFFC";
end if;
if pc = 14248 then
	inst <= x"82000844";
end if;
if pc = 14252 then
	inst <= x"07DC0018";
end if;
if pc = 14256 then
	inst <= x"C85C0008";
end if;
if pc = 14260 then
	inst <= x"48242000";
end if;
if pc = 14264 then
	inst <= x"C03C0000";
end if;
if pc = 14268 then
	inst <= x"CC220000";
end if;
if pc = 14272 then
	inst <= x"02200001";
end if;
if pc = 14276 then
	inst <= x"C1FDFFFC";
end if;
if pc = 14280 then
	inst <= x"02600000";
end if;
if pc = 14284 then
	inst <= x"02800001";
end if;
if pc = 14288 then
	inst <= x"02A00002";
end if;
if pc = 14292 then
	inst <= x"CC3C0010";
end if;
if pc = 14296 then
	inst <= x"CC7C0018";
end if;
if pc = 14300 then
	inst <= x"CC5C0020";
end if;
if pc = 14304 then
	inst <= x"C45C0028";
end if;
if pc = 14308 then
	inst <= x"C43C002C";
end if;
if pc = 14312 then
	inst <= x"C17DFFFC";
end if;
if pc = 14316 then
	inst <= x"03DC0038";
end if;
if pc = 14320 then
	inst <= x"037E000C";
end if;
if pc = 14324 then
	inst <= x"C57DFFFC";
end if;
if pc = 14328 then
	inst <= x"8200317C";
end if;
if pc = 14332 then
	inst <= x"07DC0038";
end if;
if pc = 14336 then
	inst <= x"8220380C";
end if;
if pc = 14340 then
	inst <= x"02200001";
end if;
if pc = 14344 then
	inst <= x"C1FDFFFC";
end if;
if pc = 14348 then
	inst <= x"02600001";
end if;
if pc = 14352 then
	inst <= x"02800002";
end if;
if pc = 14356 then
	inst <= x"02A00000";
end if;
if pc = 14360 then
	inst <= x"C83C0020";
end if;
if pc = 14364 then
	inst <= x"C85C0018";
end if;
if pc = 14368 then
	inst <= x"C87C0010";
end if;
if pc = 14372 then
	inst <= x"C03C002C";
end if;
if pc = 14376 then
	inst <= x"C05C0028";
end if;
if pc = 14380 then
	inst <= x"C17DFFFC";
end if;
if pc = 14384 then
	inst <= x"03DC0038";
end if;
if pc = 14388 then
	inst <= x"037E000C";
end if;
if pc = 14392 then
	inst <= x"C57DFFFC";
end if;
if pc = 14396 then
	inst <= x"8200317C";
end if;
if pc = 14400 then
	inst <= x"07DC0038";
end if;
if pc = 14404 then
	inst <= x"82203850";
end if;
if pc = 14408 then
	inst <= x"02200002";
end if;
if pc = 14412 then
	inst <= x"C1FDFFFC";
end if;
if pc = 14416 then
	inst <= x"02600002";
end if;
if pc = 14420 then
	inst <= x"02800000";
end if;
if pc = 14424 then
	inst <= x"02A00001";
end if;
if pc = 14428 then
	inst <= x"C83C0018";
end if;
if pc = 14432 then
	inst <= x"C85C0010";
end if;
if pc = 14436 then
	inst <= x"C87C0020";
end if;
if pc = 14440 then
	inst <= x"C03C002C";
end if;
if pc = 14444 then
	inst <= x"C05C0028";
end if;
if pc = 14448 then
	inst <= x"C17DFFFC";
end if;
if pc = 14452 then
	inst <= x"03DC0038";
end if;
if pc = 14456 then
	inst <= x"037E000C";
end if;
if pc = 14460 then
	inst <= x"C57DFFFC";
end if;
if pc = 14464 then
	inst <= x"8200317C";
end if;
if pc = 14468 then
	inst <= x"07DC0038";
end if;
if pc = 14472 then
	inst <= x"82203894";
end if;
if pc = 14476 then
	inst <= x"02200003";
end if;
if pc = 14480 then
	inst <= x"C1FDFFFC";
end if;
if pc = 14484 then
	inst <= x"02200000";
end if;
if pc = 14488 then
	inst <= x"C1FDFFFC";
end if;
if pc = 14492 then
	inst <= x"C8860000";
end if;
if pc = 14496 then
	inst <= x"44882000";
end if;
if pc = 14500 then
	inst <= x"C8A60004";
end if;
if pc = 14504 then
	inst <= x"4888A000";
end if;
if pc = 14508 then
	inst <= x"C8A40004";
end if;
if pc = 14512 then
	inst <= x"48A8A000";
end if;
if pc = 14516 then
	inst <= x"40AA4000";
end if;
if pc = 14520 then
	inst <= x"8EA038C0";
end if;
if pc = 14524 then
	inst <= x"820038C4";
end if;
if pc = 14528 then
	inst <= x"44A0A000";
end if;
if pc = 14532 then
	inst <= x"C0820010";
end if;
if pc = 14536 then
	inst <= x"C8C80004";
end if;
if pc = 14540 then
	inst <= x"8EAC38D8";
end if;
if pc = 14544 then
	inst <= x"02800000";
end if;
if pc = 14548 then
	inst <= x"82003918";
end if;
if pc = 14552 then
	inst <= x"C8A40008";
end if;
if pc = 14556 then
	inst <= x"48A8A000";
end if;
if pc = 14560 then
	inst <= x"40AA6000";
end if;
if pc = 14564 then
	inst <= x"8EA038EC";
end if;
if pc = 14568 then
	inst <= x"820038F0";
end if;
if pc = 14572 then
	inst <= x"44A0A000";
end if;
if pc = 14576 then
	inst <= x"C0820010";
end if;
if pc = 14580 then
	inst <= x"C8C80008";
end if;
if pc = 14584 then
	inst <= x"8EAC3904";
end if;
if pc = 14588 then
	inst <= x"02800000";
end if;
if pc = 14592 then
	inst <= x"82003918";
end if;
if pc = 14596 then
	inst <= x"C8A60004";
end if;
if pc = 14600 then
	inst <= x"8AA03914";
end if;
if pc = 14604 then
	inst <= x"02800001";
end if;
if pc = 14608 then
	inst <= x"82003918";
end if;
if pc = 14612 then
	inst <= x"02800000";
end if;
if pc = 14616 then
	inst <= x"8280392C";
end if;
if pc = 14620 then
	inst <= x"022002AC";
end if;
if pc = 14624 then
	inst <= x"CC820000";
end if;
if pc = 14628 then
	inst <= x"02200001";
end if;
if pc = 14632 then
	inst <= x"C1FDFFFC";
end if;
if pc = 14636 then
	inst <= x"C8860008";
end if;
if pc = 14640 then
	inst <= x"44884000";
end if;
if pc = 14644 then
	inst <= x"C8A6000C";
end if;
if pc = 14648 then
	inst <= x"4888A000";
end if;
if pc = 14652 then
	inst <= x"C8A40000";
end if;
if pc = 14656 then
	inst <= x"48A8A000";
end if;
if pc = 14660 then
	inst <= x"40AA2000";
end if;
if pc = 14664 then
	inst <= x"8EA03950";
end if;
if pc = 14668 then
	inst <= x"82003954";
end if;
if pc = 14672 then
	inst <= x"44A0A000";
end if;
if pc = 14676 then
	inst <= x"C0820010";
end if;
if pc = 14680 then
	inst <= x"C8C80000";
end if;
if pc = 14684 then
	inst <= x"8EAC3968";
end if;
if pc = 14688 then
	inst <= x"02800000";
end if;
if pc = 14692 then
	inst <= x"820039A8";
end if;
if pc = 14696 then
	inst <= x"C8A40008";
end if;
if pc = 14700 then
	inst <= x"48A8A000";
end if;
if pc = 14704 then
	inst <= x"40AA6000";
end if;
if pc = 14708 then
	inst <= x"8EA0397C";
end if;
if pc = 14712 then
	inst <= x"82003980";
end if;
if pc = 14716 then
	inst <= x"44A0A000";
end if;
if pc = 14720 then
	inst <= x"C0820010";
end if;
if pc = 14724 then
	inst <= x"C8C80008";
end if;
if pc = 14728 then
	inst <= x"8EAC3994";
end if;
if pc = 14732 then
	inst <= x"02800000";
end if;
if pc = 14736 then
	inst <= x"820039A8";
end if;
if pc = 14740 then
	inst <= x"C8A6000C";
end if;
if pc = 14744 then
	inst <= x"8AA039A4";
end if;
if pc = 14748 then
	inst <= x"02800001";
end if;
if pc = 14752 then
	inst <= x"820039A8";
end if;
if pc = 14756 then
	inst <= x"02800000";
end if;
if pc = 14760 then
	inst <= x"828039BC";
end if;
if pc = 14764 then
	inst <= x"022002AC";
end if;
if pc = 14768 then
	inst <= x"CC820000";
end if;
if pc = 14772 then
	inst <= x"02200002";
end if;
if pc = 14776 then
	inst <= x"C1FDFFFC";
end if;
if pc = 14780 then
	inst <= x"C8860010";
end if;
if pc = 14784 then
	inst <= x"44686000";
end if;
if pc = 14788 then
	inst <= x"C8860014";
end if;
if pc = 14792 then
	inst <= x"48668000";
end if;
if pc = 14796 then
	inst <= x"C8840000";
end if;
if pc = 14800 then
	inst <= x"48868000";
end if;
if pc = 14804 then
	inst <= x"40282000";
end if;
if pc = 14808 then
	inst <= x"8E2039E0";
end if;
if pc = 14812 then
	inst <= x"820039E4";
end if;
if pc = 14816 then
	inst <= x"44202000";
end if;
if pc = 14820 then
	inst <= x"C0820010";
end if;
if pc = 14824 then
	inst <= x"C8880000";
end if;
if pc = 14828 then
	inst <= x"8E2839F8";
end if;
if pc = 14832 then
	inst <= x"02200000";
end if;
if pc = 14836 then
	inst <= x"82003A38";
end if;
if pc = 14840 then
	inst <= x"C8240004";
end if;
if pc = 14844 then
	inst <= x"48262000";
end if;
if pc = 14848 then
	inst <= x"40224000";
end if;
if pc = 14852 then
	inst <= x"8E203A0C";
end if;
if pc = 14856 then
	inst <= x"82003A10";
end if;
if pc = 14860 then
	inst <= x"44202000";
end if;
if pc = 14864 then
	inst <= x"C0220010";
end if;
if pc = 14868 then
	inst <= x"C8420004";
end if;
if pc = 14872 then
	inst <= x"8E243A24";
end if;
if pc = 14876 then
	inst <= x"02200000";
end if;
if pc = 14880 then
	inst <= x"82003A38";
end if;
if pc = 14884 then
	inst <= x"C8260014";
end if;
if pc = 14888 then
	inst <= x"8A203A34";
end if;
if pc = 14892 then
	inst <= x"02200001";
end if;
if pc = 14896 then
	inst <= x"82003A38";
end if;
if pc = 14900 then
	inst <= x"02200000";
end if;
if pc = 14904 then
	inst <= x"82203A4C";
end if;
if pc = 14908 then
	inst <= x"022002AC";
end if;
if pc = 14912 then
	inst <= x"CC620000";
end if;
if pc = 14916 then
	inst <= x"02200003";
end if;
if pc = 14920 then
	inst <= x"C1FDFFFC";
end if;
if pc = 14924 then
	inst <= x"02200000";
end if;
if pc = 14928 then
	inst <= x"C1FDFFFC";
end if;
if pc = 14932 then
	inst <= x"C8840000";
end if;
if pc = 14936 then
	inst <= x"8A803BCC";
end if;
if pc = 14940 then
	inst <= x"C8A40004";
end if;
if pc = 14944 then
	inst <= x"48AA2000";
end if;
if pc = 14948 then
	inst <= x"C8C40008";
end if;
if pc = 14952 then
	inst <= x"48CC4000";
end if;
if pc = 14956 then
	inst <= x"40AAC000";
end if;
if pc = 14960 then
	inst <= x"C8C4000C";
end if;
if pc = 14964 then
	inst <= x"48CC6000";
end if;
if pc = 14968 then
	inst <= x"40AAC000";
end if;
if pc = 14972 then
	inst <= x"48C22000";
end if;
if pc = 14976 then
	inst <= x"C0620010";
end if;
if pc = 14980 then
	inst <= x"C8E60000";
end if;
if pc = 14984 then
	inst <= x"48CCE000";
end if;
if pc = 14988 then
	inst <= x"48E44000";
end if;
if pc = 14992 then
	inst <= x"C0620010";
end if;
if pc = 14996 then
	inst <= x"C9060004";
end if;
if pc = 15000 then
	inst <= x"48EF0000";
end if;
if pc = 15004 then
	inst <= x"40CCE000";
end if;
if pc = 15008 then
	inst <= x"48E66000";
end if;
if pc = 15012 then
	inst <= x"C0620010";
end if;
if pc = 15016 then
	inst <= x"C9060008";
end if;
if pc = 15020 then
	inst <= x"48EF0000";
end if;
if pc = 15024 then
	inst <= x"40CCE000";
end if;
if pc = 15028 then
	inst <= x"C062000C";
end if;
if pc = 15032 then
	inst <= x"82603AFC";
end if;
if pc = 15036 then
	inst <= x"48E46000";
end if;
if pc = 15040 then
	inst <= x"C0620024";
end if;
if pc = 15044 then
	inst <= x"C9060000";
end if;
if pc = 15048 then
	inst <= x"48EF0000";
end if;
if pc = 15052 then
	inst <= x"40CCE000";
end if;
if pc = 15056 then
	inst <= x"48662000";
end if;
if pc = 15060 then
	inst <= x"C0620024";
end if;
if pc = 15064 then
	inst <= x"C8E60004";
end if;
if pc = 15068 then
	inst <= x"4866E000";
end if;
if pc = 15072 then
	inst <= x"406C6000";
end if;
if pc = 15076 then
	inst <= x"48224000";
end if;
if pc = 15080 then
	inst <= x"C0620024";
end if;
if pc = 15084 then
	inst <= x"C8460008";
end if;
if pc = 15088 then
	inst <= x"48224000";
end if;
if pc = 15092 then
	inst <= x"40262000";
end if;
if pc = 15096 then
	inst <= x"82003B00";
end if;
if pc = 15100 then
	inst <= x"4020C000";
end if;
if pc = 15104 then
	inst <= x"C0620004";
end if;
if pc = 15108 then
	inst <= x"02800003";
end if;
if pc = 15112 then
	inst <= x"82683B10";
end if;
if pc = 15116 then
	inst <= x"82003B18";
end if;
if pc = 15120 then
	inst <= x"C84000A8";
end if;
if pc = 15124 then
	inst <= x"44224000";
end if;
if pc = 15128 then
	inst <= x"484AA000";
end if;
if pc = 15132 then
	inst <= x"48282000";
end if;
if pc = 15136 then
	inst <= x"44242000";
end if;
if pc = 15140 then
	inst <= x"8E023B30";
end if;
if pc = 15144 then
	inst <= x"02200000";
end if;
if pc = 15148 then
	inst <= x"C1FDFFFC";
end if;
if pc = 15152 then
	inst <= x"C0220018";
end if;
if pc = 15156 then
	inst <= x"82203B80";
end if;
if pc = 15160 then
	inst <= x"022002AC";
end if;
if pc = 15164 then
	inst <= x"C43C0000";
end if;
if pc = 15168 then
	inst <= x"C45C0004";
end if;
if pc = 15172 then
	inst <= x"CCBC0008";
end if;
if pc = 15176 then
	inst <= x"C17DFFFC";
end if;
if pc = 15180 then
	inst <= x"03DC0018";
end if;
if pc = 15184 then
	inst <= x"037E000C";
end if;
if pc = 15188 then
	inst <= x"C57DFFFC";
end if;
if pc = 15192 then
	inst <= x"8200083C";
end if;
if pc = 15196 then
	inst <= x"07DC0018";
end if;
if pc = 15200 then
	inst <= x"C85C0008";
end if;
if pc = 15204 then
	inst <= x"40242000";
end if;
if pc = 15208 then
	inst <= x"C03C0004";
end if;
if pc = 15212 then
	inst <= x"C8420010";
end if;
if pc = 15216 then
	inst <= x"48224000";
end if;
if pc = 15220 then
	inst <= x"C03C0000";
end if;
if pc = 15224 then
	inst <= x"CC220000";
end if;
if pc = 15228 then
	inst <= x"82003BC4";
end if;
if pc = 15232 then
	inst <= x"022002AC";
end if;
if pc = 15236 then
	inst <= x"C43C0010";
end if;
if pc = 15240 then
	inst <= x"C45C0004";
end if;
if pc = 15244 then
	inst <= x"CCBC0008";
end if;
if pc = 15248 then
	inst <= x"C17DFFFC";
end if;
if pc = 15252 then
	inst <= x"03DC001C";
end if;
if pc = 15256 then
	inst <= x"037E000C";
end if;
if pc = 15260 then
	inst <= x"C57DFFFC";
end if;
if pc = 15264 then
	inst <= x"8200083C";
end if;
if pc = 15268 then
	inst <= x"07DC001C";
end if;
if pc = 15272 then
	inst <= x"C85C0008";
end if;
if pc = 15276 then
	inst <= x"44242000";
end if;
if pc = 15280 then
	inst <= x"C03C0004";
end if;
if pc = 15284 then
	inst <= x"C8420010";
end if;
if pc = 15288 then
	inst <= x"48224000";
end if;
if pc = 15292 then
	inst <= x"C03C0010";
end if;
if pc = 15296 then
	inst <= x"CC220000";
end if;
if pc = 15300 then
	inst <= x"02200001";
end if;
if pc = 15304 then
	inst <= x"C1FDFFFC";
end if;
if pc = 15308 then
	inst <= x"02200000";
end if;
if pc = 15312 then
	inst <= x"C1FDFFFC";
end if;
if pc = 15316 then
	inst <= x"C8840000";
end if;
if pc = 15320 then
	inst <= x"8A803CBC";
end if;
if pc = 15324 then
	inst <= x"C8A40004";
end if;
if pc = 15328 then
	inst <= x"482A2000";
end if;
if pc = 15332 then
	inst <= x"C8A40008";
end if;
if pc = 15336 then
	inst <= x"484A4000";
end if;
if pc = 15340 then
	inst <= x"40224000";
end if;
if pc = 15344 then
	inst <= x"C844000C";
end if;
if pc = 15348 then
	inst <= x"48446000";
end if;
if pc = 15352 then
	inst <= x"40224000";
end if;
if pc = 15356 then
	inst <= x"C846000C";
end if;
if pc = 15360 then
	inst <= x"48622000";
end if;
if pc = 15364 then
	inst <= x"48484000";
end if;
if pc = 15368 then
	inst <= x"44464000";
end if;
if pc = 15372 then
	inst <= x"8E043C18";
end if;
if pc = 15376 then
	inst <= x"02200000";
end if;
if pc = 15380 then
	inst <= x"C1FDFFFC";
end if;
if pc = 15384 then
	inst <= x"C0220018";
end if;
if pc = 15388 then
	inst <= x"82203C6C";
end if;
if pc = 15392 then
	inst <= x"022002AC";
end if;
if pc = 15396 then
	inst <= x"C43C0000";
end if;
if pc = 15400 then
	inst <= x"C45C0004";
end if;
if pc = 15404 then
	inst <= x"CC3C0008";
end if;
if pc = 15408 then
	inst <= x"C17DFFFC";
end if;
if pc = 15412 then
	inst <= x"40204000";
end if;
if pc = 15416 then
	inst <= x"03DC0018";
end if;
if pc = 15420 then
	inst <= x"037E000C";
end if;
if pc = 15424 then
	inst <= x"C57DFFFC";
end if;
if pc = 15428 then
	inst <= x"8200083C";
end if;
if pc = 15432 then
	inst <= x"07DC0018";
end if;
if pc = 15436 then
	inst <= x"C85C0008";
end if;
if pc = 15440 then
	inst <= x"40242000";
end if;
if pc = 15444 then
	inst <= x"C03C0004";
end if;
if pc = 15448 then
	inst <= x"C8420010";
end if;
if pc = 15452 then
	inst <= x"48224000";
end if;
if pc = 15456 then
	inst <= x"C03C0000";
end if;
if pc = 15460 then
	inst <= x"CC220000";
end if;
if pc = 15464 then
	inst <= x"82003CB4";
end if;
if pc = 15468 then
	inst <= x"022002AC";
end if;
if pc = 15472 then
	inst <= x"C43C0010";
end if;
if pc = 15476 then
	inst <= x"C45C0004";
end if;
if pc = 15480 then
	inst <= x"CC3C0008";
end if;
if pc = 15484 then
	inst <= x"C17DFFFC";
end if;
if pc = 15488 then
	inst <= x"40204000";
end if;
if pc = 15492 then
	inst <= x"03DC001C";
end if;
if pc = 15496 then
	inst <= x"037E000C";
end if;
if pc = 15500 then
	inst <= x"C57DFFFC";
end if;
if pc = 15504 then
	inst <= x"8200083C";
end if;
if pc = 15508 then
	inst <= x"07DC001C";
end if;
if pc = 15512 then
	inst <= x"C85C0008";
end if;
if pc = 15516 then
	inst <= x"44242000";
end if;
if pc = 15520 then
	inst <= x"C03C0004";
end if;
if pc = 15524 then
	inst <= x"C8420010";
end if;
if pc = 15528 then
	inst <= x"48224000";
end if;
if pc = 15532 then
	inst <= x"C03C0010";
end if;
if pc = 15536 then
	inst <= x"CC220000";
end if;
if pc = 15540 then
	inst <= x"02200001";
end if;
if pc = 15544 then
	inst <= x"C1FDFFFC";
end if;
if pc = 15548 then
	inst <= x"02200000";
end if;
if pc = 15552 then
	inst <= x"C1FDFFFC";
end if;
if pc = 15556 then
	inst <= x"02600006";
end if;
if pc = 15560 then
	inst <= x"40200000";
end if;
if pc = 15564 then
	inst <= x"C45C0000";
end if;
if pc = 15568 then
	inst <= x"C43C0004";
end if;
if pc = 15572 then
	inst <= x"C17DFFFC";
end if;
if pc = 15576 then
	inst <= x"00260000";
end if;
if pc = 15580 then
	inst <= x"03DC0010";
end if;
if pc = 15584 then
	inst <= x"037E000C";
end if;
if pc = 15588 then
	inst <= x"C57DFFFC";
end if;
if pc = 15592 then
	inst <= x"8200081C";
end if;
if pc = 15596 then
	inst <= x"07DC0010";
end if;
if pc = 15600 then
	inst <= x"C05C0004";
end if;
if pc = 15604 then
	inst <= x"C8240000";
end if;
if pc = 15608 then
	inst <= x"8A203D78";
end if;
if pc = 15612 then
	inst <= x"C07C0000";
end if;
if pc = 15616 then
	inst <= x"C0860018";
end if;
if pc = 15620 then
	inst <= x"C8240000";
end if;
if pc = 15624 then
	inst <= x"8E203D14";
end if;
if pc = 15628 then
	inst <= x"02A00000";
end if;
if pc = 15632 then
	inst <= x"82003D18";
end if;
if pc = 15636 then
	inst <= x"02A00001";
end if;
if pc = 15640 then
	inst <= x"82803D30";
end if;
if pc = 15644 then
	inst <= x"8E203D28";
end if;
if pc = 15648 then
	inst <= x"02800001";
end if;
if pc = 15652 then
	inst <= x"82003D2C";
end if;
if pc = 15656 then
	inst <= x"02800000";
end if;
if pc = 15660 then
	inst <= x"82003D34";
end if;
if pc = 15664 then
	inst <= x"008A0000";
end if;
if pc = 15668 then
	inst <= x"C0A60010";
end if;
if pc = 15672 then
	inst <= x"C82A0000";
end if;
if pc = 15676 then
	inst <= x"82803D44";
end if;
if pc = 15680 then
	inst <= x"82003D48";
end if;
if pc = 15684 then
	inst <= x"44202000";
end if;
if pc = 15688 then
	inst <= x"CC220000";
end if;
if pc = 15692 then
	inst <= x"C8240000";
end if;
if pc = 15696 then
	inst <= x"C43C0008";
end if;
if pc = 15700 then
	inst <= x"C17DFFFC";
end if;
if pc = 15704 then
	inst <= x"03DC0014";
end if;
if pc = 15708 then
	inst <= x"037E000C";
end if;
if pc = 15712 then
	inst <= x"C57DFFFC";
end if;
if pc = 15716 then
	inst <= x"82000844";
end if;
if pc = 15720 then
	inst <= x"07DC0014";
end if;
if pc = 15724 then
	inst <= x"C03C0008";
end if;
if pc = 15728 then
	inst <= x"CC220004";
end if;
if pc = 15732 then
	inst <= x"82003D7C";
end if;
if pc = 15736 then
	inst <= x"CC020004";
end if;
if pc = 15740 then
	inst <= x"C05C0004";
end if;
if pc = 15744 then
	inst <= x"C8240004";
end if;
if pc = 15748 then
	inst <= x"8A203E04";
end if;
if pc = 15752 then
	inst <= x"C07C0000";
end if;
if pc = 15756 then
	inst <= x"C0860018";
end if;
if pc = 15760 then
	inst <= x"C8240004";
end if;
if pc = 15764 then
	inst <= x"8E203DA0";
end if;
if pc = 15768 then
	inst <= x"02A00000";
end if;
if pc = 15772 then
	inst <= x"82003DA4";
end if;
if pc = 15776 then
	inst <= x"02A00001";
end if;
if pc = 15780 then
	inst <= x"82803DBC";
end if;
if pc = 15784 then
	inst <= x"8E203DB4";
end if;
if pc = 15788 then
	inst <= x"02800001";
end if;
if pc = 15792 then
	inst <= x"82003DB8";
end if;
if pc = 15796 then
	inst <= x"02800000";
end if;
if pc = 15800 then
	inst <= x"82003DC0";
end if;
if pc = 15804 then
	inst <= x"008A0000";
end if;
if pc = 15808 then
	inst <= x"C0A60010";
end if;
if pc = 15812 then
	inst <= x"C82A0004";
end if;
if pc = 15816 then
	inst <= x"82803DD0";
end if;
if pc = 15820 then
	inst <= x"82003DD4";
end if;
if pc = 15824 then
	inst <= x"44202000";
end if;
if pc = 15828 then
	inst <= x"CC220008";
end if;
if pc = 15832 then
	inst <= x"C8240004";
end if;
if pc = 15836 then
	inst <= x"C43C0008";
end if;
if pc = 15840 then
	inst <= x"C17DFFFC";
end if;
if pc = 15844 then
	inst <= x"03DC0014";
end if;
if pc = 15848 then
	inst <= x"037E000C";
end if;
if pc = 15852 then
	inst <= x"C57DFFFC";
end if;
if pc = 15856 then
	inst <= x"82000844";
end if;
if pc = 15860 then
	inst <= x"07DC0014";
end if;
if pc = 15864 then
	inst <= x"C03C0008";
end if;
if pc = 15868 then
	inst <= x"CC22000C";
end if;
if pc = 15872 then
	inst <= x"82003E08";
end if;
if pc = 15876 then
	inst <= x"CC02000C";
end if;
if pc = 15880 then
	inst <= x"C05C0004";
end if;
if pc = 15884 then
	inst <= x"C8240008";
end if;
if pc = 15888 then
	inst <= x"8A203E90";
end if;
if pc = 15892 then
	inst <= x"C07C0000";
end if;
if pc = 15896 then
	inst <= x"C0860018";
end if;
if pc = 15900 then
	inst <= x"C8240008";
end if;
if pc = 15904 then
	inst <= x"8E203E2C";
end if;
if pc = 15908 then
	inst <= x"02A00000";
end if;
if pc = 15912 then
	inst <= x"82003E30";
end if;
if pc = 15916 then
	inst <= x"02A00001";
end if;
if pc = 15920 then
	inst <= x"82803E48";
end if;
if pc = 15924 then
	inst <= x"8E203E40";
end if;
if pc = 15928 then
	inst <= x"02800001";
end if;
if pc = 15932 then
	inst <= x"82003E44";
end if;
if pc = 15936 then
	inst <= x"02800000";
end if;
if pc = 15940 then
	inst <= x"82003E4C";
end if;
if pc = 15944 then
	inst <= x"008A0000";
end if;
if pc = 15948 then
	inst <= x"C0660010";
end if;
if pc = 15952 then
	inst <= x"C8260008";
end if;
if pc = 15956 then
	inst <= x"82803E5C";
end if;
if pc = 15960 then
	inst <= x"82003E60";
end if;
if pc = 15964 then
	inst <= x"44202000";
end if;
if pc = 15968 then
	inst <= x"CC220010";
end if;
if pc = 15972 then
	inst <= x"C8240008";
end if;
if pc = 15976 then
	inst <= x"C43C0008";
end if;
if pc = 15980 then
	inst <= x"C17DFFFC";
end if;
if pc = 15984 then
	inst <= x"03DC0014";
end if;
if pc = 15988 then
	inst <= x"037E000C";
end if;
if pc = 15992 then
	inst <= x"C57DFFFC";
end if;
if pc = 15996 then
	inst <= x"82000844";
end if;
if pc = 16000 then
	inst <= x"07DC0014";
end if;
if pc = 16004 then
	inst <= x"C03C0008";
end if;
if pc = 16008 then
	inst <= x"CC220014";
end if;
if pc = 16012 then
	inst <= x"82003E94";
end if;
if pc = 16016 then
	inst <= x"CC020014";
end if;
if pc = 16020 then
	inst <= x"C1FDFFFC";
end if;
if pc = 16024 then
	inst <= x"02600004";
end if;
if pc = 16028 then
	inst <= x"40200000";
end if;
if pc = 16032 then
	inst <= x"C45C0000";
end if;
if pc = 16036 then
	inst <= x"C43C0004";
end if;
if pc = 16040 then
	inst <= x"C17DFFFC";
end if;
if pc = 16044 then
	inst <= x"00260000";
end if;
if pc = 16048 then
	inst <= x"03DC0010";
end if;
if pc = 16052 then
	inst <= x"037E000C";
end if;
if pc = 16056 then
	inst <= x"C57DFFFC";
end if;
if pc = 16060 then
	inst <= x"8200081C";
end if;
if pc = 16064 then
	inst <= x"07DC0010";
end if;
if pc = 16068 then
	inst <= x"C05C0004";
end if;
if pc = 16072 then
	inst <= x"C8240000";
end if;
if pc = 16076 then
	inst <= x"C07C0000";
end if;
if pc = 16080 then
	inst <= x"C0860010";
end if;
if pc = 16084 then
	inst <= x"C8480000";
end if;
if pc = 16088 then
	inst <= x"48224000";
end if;
if pc = 16092 then
	inst <= x"C8440004";
end if;
if pc = 16096 then
	inst <= x"C0860010";
end if;
if pc = 16100 then
	inst <= x"C8680004";
end if;
if pc = 16104 then
	inst <= x"48446000";
end if;
if pc = 16108 then
	inst <= x"40224000";
end if;
if pc = 16112 then
	inst <= x"C8440008";
end if;
if pc = 16116 then
	inst <= x"C0460010";
end if;
if pc = 16120 then
	inst <= x"C8640008";
end if;
if pc = 16124 then
	inst <= x"48446000";
end if;
if pc = 16128 then
	inst <= x"40224000";
end if;
if pc = 16132 then
	inst <= x"8E023F10";
end if;
if pc = 16136 then
	inst <= x"CC020000";
end if;
if pc = 16140 then
	inst <= x"82004008";
end if;
if pc = 16144 then
	inst <= x"CC3C0008";
end if;
if pc = 16148 then
	inst <= x"C43C0010";
end if;
if pc = 16152 then
	inst <= x"C17DFFFC";
end if;
if pc = 16156 then
	inst <= x"03DC001C";
end if;
if pc = 16160 then
	inst <= x"037E000C";
end if;
if pc = 16164 then
	inst <= x"C57DFFFC";
end if;
if pc = 16168 then
	inst <= x"82000844";
end if;
if pc = 16172 then
	inst <= x"07DC001C";
end if;
if pc = 16176 then
	inst <= x"44202000";
end if;
if pc = 16180 then
	inst <= x"C03C0010";
end if;
if pc = 16184 then
	inst <= x"CC220000";
end if;
if pc = 16188 then
	inst <= x"C05C0000";
end if;
if pc = 16192 then
	inst <= x"C0640010";
end if;
if pc = 16196 then
	inst <= x"C8260000";
end if;
if pc = 16200 then
	inst <= x"C85C0008";
end if;
if pc = 16204 then
	inst <= x"CC3C0018";
end if;
if pc = 16208 then
	inst <= x"C17DFFFC";
end if;
if pc = 16212 then
	inst <= x"40204000";
end if;
if pc = 16216 then
	inst <= x"03DC0028";
end if;
if pc = 16220 then
	inst <= x"037E000C";
end if;
if pc = 16224 then
	inst <= x"C57DFFFC";
end if;
if pc = 16228 then
	inst <= x"82000844";
end if;
if pc = 16232 then
	inst <= x"07DC0028";
end if;
if pc = 16236 then
	inst <= x"C85C0018";
end if;
if pc = 16240 then
	inst <= x"48242000";
end if;
if pc = 16244 then
	inst <= x"44202000";
end if;
if pc = 16248 then
	inst <= x"C03C0010";
end if;
if pc = 16252 then
	inst <= x"CC220004";
end if;
if pc = 16256 then
	inst <= x"C05C0000";
end if;
if pc = 16260 then
	inst <= x"C0640010";
end if;
if pc = 16264 then
	inst <= x"C8260004";
end if;
if pc = 16268 then
	inst <= x"C85C0008";
end if;
if pc = 16272 then
	inst <= x"CC3C0020";
end if;
if pc = 16276 then
	inst <= x"C17DFFFC";
end if;
if pc = 16280 then
	inst <= x"40204000";
end if;
if pc = 16284 then
	inst <= x"03DC0030";
end if;
if pc = 16288 then
	inst <= x"037E000C";
end if;
if pc = 16292 then
	inst <= x"C57DFFFC";
end if;
if pc = 16296 then
	inst <= x"82000844";
end if;
if pc = 16300 then
	inst <= x"07DC0030";
end if;
if pc = 16304 then
	inst <= x"C85C0020";
end if;
if pc = 16308 then
	inst <= x"48242000";
end if;
if pc = 16312 then
	inst <= x"44202000";
end if;
if pc = 16316 then
	inst <= x"C03C0010";
end if;
if pc = 16320 then
	inst <= x"CC220008";
end if;
if pc = 16324 then
	inst <= x"C05C0000";
end if;
if pc = 16328 then
	inst <= x"C0440010";
end if;
if pc = 16332 then
	inst <= x"C8240008";
end if;
if pc = 16336 then
	inst <= x"C85C0008";
end if;
if pc = 16340 then
	inst <= x"CC3C0028";
end if;
if pc = 16344 then
	inst <= x"C17DFFFC";
end if;
if pc = 16348 then
	inst <= x"40204000";
end if;
if pc = 16352 then
	inst <= x"03DC0038";
end if;
if pc = 16356 then
	inst <= x"037E000C";
end if;
if pc = 16360 then
	inst <= x"C57DFFFC";
end if;
if pc = 16364 then
	inst <= x"82000844";
end if;
if pc = 16368 then
	inst <= x"07DC0038";
end if;
if pc = 16372 then
	inst <= x"C85C0028";
end if;
if pc = 16376 then
	inst <= x"48242000";
end if;
if pc = 16380 then
	inst <= x"44202000";
end if;
if pc = 16384 then
	inst <= x"C03C0010";
end if;
if pc = 16388 then
	inst <= x"CC22000C";
end if;
if pc = 16392 then
	inst <= x"C1FDFFFC";
end if;
if pc = 16396 then
	inst <= x"02600005";
end if;
if pc = 16400 then
	inst <= x"40200000";
end if;
if pc = 16404 then
	inst <= x"C45C0000";
end if;
if pc = 16408 then
	inst <= x"C43C0004";
end if;
if pc = 16412 then
	inst <= x"C17DFFFC";
end if;
if pc = 16416 then
	inst <= x"00260000";
end if;
if pc = 16420 then
	inst <= x"03DC0010";
end if;
if pc = 16424 then
	inst <= x"037E000C";
end if;
if pc = 16428 then
	inst <= x"C57DFFFC";
end if;
if pc = 16432 then
	inst <= x"8200081C";
end if;
if pc = 16436 then
	inst <= x"07DC0010";
end if;
if pc = 16440 then
	inst <= x"C05C0004";
end if;
if pc = 16444 then
	inst <= x"C8240000";
end if;
if pc = 16448 then
	inst <= x"C8440004";
end if;
if pc = 16452 then
	inst <= x"C8640008";
end if;
if pc = 16456 then
	inst <= x"48822000";
end if;
if pc = 16460 then
	inst <= x"C07C0000";
end if;
if pc = 16464 then
	inst <= x"C0860010";
end if;
if pc = 16468 then
	inst <= x"C8A80000";
end if;
if pc = 16472 then
	inst <= x"4888A000";
end if;
if pc = 16476 then
	inst <= x"48A44000";
end if;
if pc = 16480 then
	inst <= x"C0860010";
end if;
if pc = 16484 then
	inst <= x"C8C80004";
end if;
if pc = 16488 then
	inst <= x"48AAC000";
end if;
if pc = 16492 then
	inst <= x"4088A000";
end if;
if pc = 16496 then
	inst <= x"48A66000";
end if;
if pc = 16500 then
	inst <= x"C0860010";
end if;
if pc = 16504 then
	inst <= x"C8C80008";
end if;
if pc = 16508 then
	inst <= x"48AAC000";
end if;
if pc = 16512 then
	inst <= x"4088A000";
end if;
if pc = 16516 then
	inst <= x"C086000C";
end if;
if pc = 16520 then
	inst <= x"828040CC";
end if;
if pc = 16524 then
	inst <= x"48A46000";
end if;
if pc = 16528 then
	inst <= x"C0860024";
end if;
if pc = 16532 then
	inst <= x"C8C80000";
end if;
if pc = 16536 then
	inst <= x"48AAC000";
end if;
if pc = 16540 then
	inst <= x"4088A000";
end if;
if pc = 16544 then
	inst <= x"48662000";
end if;
if pc = 16548 then
	inst <= x"C0860024";
end if;
if pc = 16552 then
	inst <= x"C8A80004";
end if;
if pc = 16556 then
	inst <= x"4866A000";
end if;
if pc = 16560 then
	inst <= x"40686000";
end if;
if pc = 16564 then
	inst <= x"48224000";
end if;
if pc = 16568 then
	inst <= x"C0860024";
end if;
if pc = 16572 then
	inst <= x"C8480008";
end if;
if pc = 16576 then
	inst <= x"48224000";
end if;
if pc = 16580 then
	inst <= x"40262000";
end if;
if pc = 16584 then
	inst <= x"820040D0";
end if;
if pc = 16588 then
	inst <= x"40208000";
end if;
if pc = 16592 then
	inst <= x"C8440000";
end if;
if pc = 16596 then
	inst <= x"C0860010";
end if;
if pc = 16600 then
	inst <= x"C8680000";
end if;
if pc = 16604 then
	inst <= x"48446000";
end if;
if pc = 16608 then
	inst <= x"44404000";
end if;
if pc = 16612 then
	inst <= x"C8640004";
end if;
if pc = 16616 then
	inst <= x"C0860010";
end if;
if pc = 16620 then
	inst <= x"C8880004";
end if;
if pc = 16624 then
	inst <= x"48668000";
end if;
if pc = 16628 then
	inst <= x"44606000";
end if;
if pc = 16632 then
	inst <= x"C8840008";
end if;
if pc = 16636 then
	inst <= x"C0860010";
end if;
if pc = 16640 then
	inst <= x"C8A80008";
end if;
if pc = 16644 then
	inst <= x"4888A000";
end if;
if pc = 16648 then
	inst <= x"44808000";
end if;
if pc = 16652 then
	inst <= x"CC220000";
end if;
if pc = 16656 then
	inst <= x"C086000C";
end if;
if pc = 16660 then
	inst <= x"CC3C0008";
end if;
if pc = 16664 then
	inst <= x"82804264";
end if;
if pc = 16668 then
	inst <= x"C8A40008";
end if;
if pc = 16672 then
	inst <= x"C0860024";
end if;
if pc = 16676 then
	inst <= x"C8C80004";
end if;
if pc = 16680 then
	inst <= x"48AAC000";
end if;
if pc = 16684 then
	inst <= x"C8C40004";
end if;
if pc = 16688 then
	inst <= x"C0860024";
end if;
if pc = 16692 then
	inst <= x"C8E80008";
end if;
if pc = 16696 then
	inst <= x"48CCE000";
end if;
if pc = 16700 then
	inst <= x"40AAC000";
end if;
if pc = 16704 then
	inst <= x"C8C00080";
end if;
if pc = 16708 then
	inst <= x"CC9C0010";
end if;
if pc = 16712 then
	inst <= x"CC7C0018";
end if;
if pc = 16716 then
	inst <= x"CCDC0020";
end if;
if pc = 16720 then
	inst <= x"C43C0028";
end if;
if pc = 16724 then
	inst <= x"CC5C0030";
end if;
if pc = 16728 then
	inst <= x"CCBC0038";
end if;
if pc = 16732 then
	inst <= x"C17DFFFC";
end if;
if pc = 16736 then
	inst <= x"4020C000";
end if;
if pc = 16740 then
	inst <= x"03DC0048";
end if;
if pc = 16744 then
	inst <= x"037E000C";
end if;
if pc = 16748 then
	inst <= x"C57DFFFC";
end if;
if pc = 16752 then
	inst <= x"82000844";
end if;
if pc = 16756 then
	inst <= x"07DC0048";
end if;
if pc = 16760 then
	inst <= x"C85C0038";
end if;
if pc = 16764 then
	inst <= x"48242000";
end if;
if pc = 16768 then
	inst <= x"C85C0030";
end if;
if pc = 16772 then
	inst <= x"44242000";
end if;
if pc = 16776 then
	inst <= x"C03C0028";
end if;
if pc = 16780 then
	inst <= x"CC220004";
end if;
if pc = 16784 then
	inst <= x"C05C0004";
end if;
if pc = 16788 then
	inst <= x"C8240008";
end if;
if pc = 16792 then
	inst <= x"C07C0000";
end if;
if pc = 16796 then
	inst <= x"C0860024";
end if;
if pc = 16800 then
	inst <= x"C8480000";
end if;
if pc = 16804 then
	inst <= x"48224000";
end if;
if pc = 16808 then
	inst <= x"C8440000";
end if;
if pc = 16812 then
	inst <= x"C0860024";
end if;
if pc = 16816 then
	inst <= x"C8680008";
end if;
if pc = 16820 then
	inst <= x"48446000";
end if;
if pc = 16824 then
	inst <= x"40224000";
end if;
if pc = 16828 then
	inst <= x"C85C0020";
end if;
if pc = 16832 then
	inst <= x"CC3C0040";
end if;
if pc = 16836 then
	inst <= x"C17DFFFC";
end if;
if pc = 16840 then
	inst <= x"40204000";
end if;
if pc = 16844 then
	inst <= x"03DC0050";
end if;
if pc = 16848 then
	inst <= x"037E000C";
end if;
if pc = 16852 then
	inst <= x"C57DFFFC";
end if;
if pc = 16856 then
	inst <= x"82000844";
end if;
if pc = 16860 then
	inst <= x"07DC0050";
end if;
if pc = 16864 then
	inst <= x"C85C0040";
end if;
if pc = 16868 then
	inst <= x"48242000";
end if;
if pc = 16872 then
	inst <= x"C85C0018";
end if;
if pc = 16876 then
	inst <= x"44242000";
end if;
if pc = 16880 then
	inst <= x"C03C0028";
end if;
if pc = 16884 then
	inst <= x"CC220008";
end if;
if pc = 16888 then
	inst <= x"C05C0004";
end if;
if pc = 16892 then
	inst <= x"C8240004";
end if;
if pc = 16896 then
	inst <= x"C07C0000";
end if;
if pc = 16900 then
	inst <= x"C0860024";
end if;
if pc = 16904 then
	inst <= x"C8480000";
end if;
if pc = 16908 then
	inst <= x"48224000";
end if;
if pc = 16912 then
	inst <= x"C8440000";
end if;
if pc = 16916 then
	inst <= x"C0460024";
end if;
if pc = 16920 then
	inst <= x"C8640004";
end if;
if pc = 16924 then
	inst <= x"48446000";
end if;
if pc = 16928 then
	inst <= x"40224000";
end if;
if pc = 16932 then
	inst <= x"C85C0020";
end if;
if pc = 16936 then
	inst <= x"CC3C0048";
end if;
if pc = 16940 then
	inst <= x"C17DFFFC";
end if;
if pc = 16944 then
	inst <= x"40204000";
end if;
if pc = 16948 then
	inst <= x"03DC0058";
end if;
if pc = 16952 then
	inst <= x"037E000C";
end if;
if pc = 16956 then
	inst <= x"C57DFFFC";
end if;
if pc = 16960 then
	inst <= x"82000844";
end if;
if pc = 16964 then
	inst <= x"07DC0058";
end if;
if pc = 16968 then
	inst <= x"C85C0048";
end if;
if pc = 16972 then
	inst <= x"48242000";
end if;
if pc = 16976 then
	inst <= x"C85C0010";
end if;
if pc = 16980 then
	inst <= x"44242000";
end if;
if pc = 16984 then
	inst <= x"C03C0028";
end if;
if pc = 16988 then
	inst <= x"CC22000C";
end if;
if pc = 16992 then
	inst <= x"82004270";
end if;
if pc = 16996 then
	inst <= x"CC420004";
end if;
if pc = 17000 then
	inst <= x"CC620008";
end if;
if pc = 17004 then
	inst <= x"CC82000C";
end if;
if pc = 17008 then
	inst <= x"C83C0008";
end if;
if pc = 17012 then
	inst <= x"8A2042A0";
end if;
if pc = 17016 then
	inst <= x"C43C0028";
end if;
if pc = 17020 then
	inst <= x"C17DFFFC";
end if;
if pc = 17024 then
	inst <= x"03DC0058";
end if;
if pc = 17028 then
	inst <= x"037E000C";
end if;
if pc = 17032 then
	inst <= x"C57DFFFC";
end if;
if pc = 17036 then
	inst <= x"82000844";
end if;
if pc = 17040 then
	inst <= x"07DC0058";
end if;
if pc = 17044 then
	inst <= x"C03C0028";
end if;
if pc = 17048 then
	inst <= x"CC220010";
end if;
if pc = 17052 then
	inst <= x"820042A0";
end if;
if pc = 17056 then
	inst <= x"C1FDFFFC";
end if;
if pc = 17060 then
	inst <= x"86404628";
end if;
if pc = 17064 then
	inst <= x"026000C8";
end if;
if pc = 17068 then
	inst <= x"22840220";
end if;
if pc = 17072 then
	inst <= x"D0868000";
end if;
if pc = 17076 then
	inst <= x"C0A20004";
end if;
if pc = 17080 then
	inst <= x"C0C20000";
end if;
if pc = 17084 then
	inst <= x"C0E80004";
end if;
if pc = 17088 then
	inst <= x"03000001";
end if;
if pc = 17092 then
	inst <= x"C43C0000";
end if;
if pc = 17096 then
	inst <= x"C47C0004";
end if;
if pc = 17100 then
	inst <= x"82F04350";
end if;
if pc = 17104 then
	inst <= x"03000002";
end if;
if pc = 17108 then
	inst <= x"82F04314";
end if;
if pc = 17112 then
	inst <= x"C4BC0008";
end if;
if pc = 17116 then
	inst <= x"C45C000C";
end if;
if pc = 17120 then
	inst <= x"C17DFFFC";
end if;
if pc = 17124 then
	inst <= x"00480000";
end if;
if pc = 17128 then
	inst <= x"002C0000";
end if;
if pc = 17132 then
	inst <= x"03DC0018";
end if;
if pc = 17136 then
	inst <= x"037E000C";
end if;
if pc = 17140 then
	inst <= x"C57DFFFC";
end if;
if pc = 17144 then
	inst <= x"8200400C";
end if;
if pc = 17148 then
	inst <= x"07DC0018";
end if;
if pc = 17152 then
	inst <= x"C05C000C";
end if;
if pc = 17156 then
	inst <= x"22640220";
end if;
if pc = 17160 then
	inst <= x"C09C0008";
end if;
if pc = 17164 then
	inst <= x"D4286000";
end if;
if pc = 17168 then
	inst <= x"8200434C";
end if;
if pc = 17172 then
	inst <= x"C4BC0008";
end if;
if pc = 17176 then
	inst <= x"C45C000C";
end if;
if pc = 17180 then
	inst <= x"C17DFFFC";
end if;
if pc = 17184 then
	inst <= x"00480000";
end if;
if pc = 17188 then
	inst <= x"002C0000";
end if;
if pc = 17192 then
	inst <= x"03DC0018";
end if;
if pc = 17196 then
	inst <= x"037E000C";
end if;
if pc = 17200 then
	inst <= x"C57DFFFC";
end if;
if pc = 17204 then
	inst <= x"82003E98";
end if;
if pc = 17208 then
	inst <= x"07DC0018";
end if;
if pc = 17212 then
	inst <= x"C05C000C";
end if;
if pc = 17216 then
	inst <= x"22640220";
end if;
if pc = 17220 then
	inst <= x"C09C0008";
end if;
if pc = 17224 then
	inst <= x"D4286000";
end if;
if pc = 17228 then
	inst <= x"82004388";
end if;
if pc = 17232 then
	inst <= x"C4BC0008";
end if;
if pc = 17236 then
	inst <= x"C45C000C";
end if;
if pc = 17240 then
	inst <= x"C17DFFFC";
end if;
if pc = 17244 then
	inst <= x"00480000";
end if;
if pc = 17248 then
	inst <= x"002C0000";
end if;
if pc = 17252 then
	inst <= x"03DC0018";
end if;
if pc = 17256 then
	inst <= x"037E000C";
end if;
if pc = 17260 then
	inst <= x"C57DFFFC";
end if;
if pc = 17264 then
	inst <= x"82003CC4";
end if;
if pc = 17268 then
	inst <= x"07DC0018";
end if;
if pc = 17272 then
	inst <= x"C05C000C";
end if;
if pc = 17276 then
	inst <= x"22640220";
end if;
if pc = 17280 then
	inst <= x"C09C0008";
end if;
if pc = 17284 then
	inst <= x"D4286000";
end if;
if pc = 17288 then
	inst <= x"06240001";
end if;
if pc = 17292 then
	inst <= x"86204624";
end if;
if pc = 17296 then
	inst <= x"22420220";
end if;
if pc = 17300 then
	inst <= x"C07C0004";
end if;
if pc = 17304 then
	inst <= x"D0464000";
end if;
if pc = 17308 then
	inst <= x"C09C0000";
end if;
if pc = 17312 then
	inst <= x"C0A80004";
end if;
if pc = 17316 then
	inst <= x"C0C80000";
end if;
if pc = 17320 then
	inst <= x"C0E40004";
end if;
if pc = 17324 then
	inst <= x"03000001";
end if;
if pc = 17328 then
	inst <= x"82F0442C";
end if;
if pc = 17332 then
	inst <= x"03000002";
end if;
if pc = 17336 then
	inst <= x"82F043F4";
end if;
if pc = 17340 then
	inst <= x"C4BC0010";
end if;
if pc = 17344 then
	inst <= x"C43C0014";
end if;
if pc = 17348 then
	inst <= x"C17DFFFC";
end if;
if pc = 17352 then
	inst <= x"002C0000";
end if;
if pc = 17356 then
	inst <= x"03DC0020";
end if;
if pc = 17360 then
	inst <= x"037E000C";
end if;
if pc = 17364 then
	inst <= x"C57DFFFC";
end if;
if pc = 17368 then
	inst <= x"8200400C";
end if;
if pc = 17372 then
	inst <= x"07DC0020";
end if;
if pc = 17376 then
	inst <= x"C05C0014";
end if;
if pc = 17380 then
	inst <= x"22640220";
end if;
if pc = 17384 then
	inst <= x"C09C0010";
end if;
if pc = 17388 then
	inst <= x"D4286000";
end if;
if pc = 17392 then
	inst <= x"82004428";
end if;
if pc = 17396 then
	inst <= x"C4BC0010";
end if;
if pc = 17400 then
	inst <= x"C43C0014";
end if;
if pc = 17404 then
	inst <= x"C17DFFFC";
end if;
if pc = 17408 then
	inst <= x"002C0000";
end if;
if pc = 17412 then
	inst <= x"03DC0020";
end if;
if pc = 17416 then
	inst <= x"037E000C";
end if;
if pc = 17420 then
	inst <= x"C57DFFFC";
end if;
if pc = 17424 then
	inst <= x"82003E98";
end if;
if pc = 17428 then
	inst <= x"07DC0020";
end if;
if pc = 17432 then
	inst <= x"C05C0014";
end if;
if pc = 17436 then
	inst <= x"22640220";
end if;
if pc = 17440 then
	inst <= x"C09C0010";
end if;
if pc = 17444 then
	inst <= x"D4286000";
end if;
if pc = 17448 then
	inst <= x"82004460";
end if;
if pc = 17452 then
	inst <= x"C4BC0010";
end if;
if pc = 17456 then
	inst <= x"C43C0014";
end if;
if pc = 17460 then
	inst <= x"C17DFFFC";
end if;
if pc = 17464 then
	inst <= x"002C0000";
end if;
if pc = 17468 then
	inst <= x"03DC0020";
end if;
if pc = 17472 then
	inst <= x"037E000C";
end if;
if pc = 17476 then
	inst <= x"C57DFFFC";
end if;
if pc = 17480 then
	inst <= x"82003CC4";
end if;
if pc = 17484 then
	inst <= x"07DC0020";
end if;
if pc = 17488 then
	inst <= x"C05C0014";
end if;
if pc = 17492 then
	inst <= x"22640220";
end if;
if pc = 17496 then
	inst <= x"C09C0010";
end if;
if pc = 17500 then
	inst <= x"D4286000";
end if;
if pc = 17504 then
	inst <= x"06240001";
end if;
if pc = 17508 then
	inst <= x"86204620";
end if;
if pc = 17512 then
	inst <= x"22420220";
end if;
if pc = 17516 then
	inst <= x"C07C0004";
end if;
if pc = 17520 then
	inst <= x"D0464000";
end if;
if pc = 17524 then
	inst <= x"C09C0000";
end if;
if pc = 17528 then
	inst <= x"C0A80004";
end if;
if pc = 17532 then
	inst <= x"C0C80000";
end if;
if pc = 17536 then
	inst <= x"C0E40004";
end if;
if pc = 17540 then
	inst <= x"03000001";
end if;
if pc = 17544 then
	inst <= x"82F04504";
end if;
if pc = 17548 then
	inst <= x"03000002";
end if;
if pc = 17552 then
	inst <= x"82F044CC";
end if;
if pc = 17556 then
	inst <= x"C4BC0018";
end if;
if pc = 17560 then
	inst <= x"C43C001C";
end if;
if pc = 17564 then
	inst <= x"C17DFFFC";
end if;
if pc = 17568 then
	inst <= x"002C0000";
end if;
if pc = 17572 then
	inst <= x"03DC0028";
end if;
if pc = 17576 then
	inst <= x"037E000C";
end if;
if pc = 17580 then
	inst <= x"C57DFFFC";
end if;
if pc = 17584 then
	inst <= x"8200400C";
end if;
if pc = 17588 then
	inst <= x"07DC0028";
end if;
if pc = 17592 then
	inst <= x"C05C001C";
end if;
if pc = 17596 then
	inst <= x"22640220";
end if;
if pc = 17600 then
	inst <= x"C09C0018";
end if;
if pc = 17604 then
	inst <= x"D4286000";
end if;
if pc = 17608 then
	inst <= x"82004500";
end if;
if pc = 17612 then
	inst <= x"C4BC0018";
end if;
if pc = 17616 then
	inst <= x"C43C001C";
end if;
if pc = 17620 then
	inst <= x"C17DFFFC";
end if;
if pc = 17624 then
	inst <= x"002C0000";
end if;
if pc = 17628 then
	inst <= x"03DC0028";
end if;
if pc = 17632 then
	inst <= x"037E000C";
end if;
if pc = 17636 then
	inst <= x"C57DFFFC";
end if;
if pc = 17640 then
	inst <= x"82003E98";
end if;
if pc = 17644 then
	inst <= x"07DC0028";
end if;
if pc = 17648 then
	inst <= x"C05C001C";
end if;
if pc = 17652 then
	inst <= x"22640220";
end if;
if pc = 17656 then
	inst <= x"C09C0018";
end if;
if pc = 17660 then
	inst <= x"D4286000";
end if;
if pc = 17664 then
	inst <= x"82004538";
end if;
if pc = 17668 then
	inst <= x"C4BC0018";
end if;
if pc = 17672 then
	inst <= x"C43C001C";
end if;
if pc = 17676 then
	inst <= x"C17DFFFC";
end if;
if pc = 17680 then
	inst <= x"002C0000";
end if;
if pc = 17684 then
	inst <= x"03DC0028";
end if;
if pc = 17688 then
	inst <= x"037E000C";
end if;
if pc = 17692 then
	inst <= x"C57DFFFC";
end if;
if pc = 17696 then
	inst <= x"82003CC4";
end if;
if pc = 17700 then
	inst <= x"07DC0028";
end if;
if pc = 17704 then
	inst <= x"C05C001C";
end if;
if pc = 17708 then
	inst <= x"22640220";
end if;
if pc = 17712 then
	inst <= x"C09C0018";
end if;
if pc = 17716 then
	inst <= x"D4286000";
end if;
if pc = 17720 then
	inst <= x"06240001";
end if;
if pc = 17724 then
	inst <= x"8620461C";
end if;
if pc = 17728 then
	inst <= x"22420220";
end if;
if pc = 17732 then
	inst <= x"C07C0004";
end if;
if pc = 17736 then
	inst <= x"D0464000";
end if;
if pc = 17740 then
	inst <= x"C07C0000";
end if;
if pc = 17744 then
	inst <= x"C0860004";
end if;
if pc = 17748 then
	inst <= x"C0A60000";
end if;
if pc = 17752 then
	inst <= x"C0C40004";
end if;
if pc = 17756 then
	inst <= x"02E00001";
end if;
if pc = 17760 then
	inst <= x"82CE45DC";
end if;
if pc = 17764 then
	inst <= x"02E00002";
end if;
if pc = 17768 then
	inst <= x"82CE45A4";
end if;
if pc = 17772 then
	inst <= x"C49C0020";
end if;
if pc = 17776 then
	inst <= x"C43C0024";
end if;
if pc = 17780 then
	inst <= x"C17DFFFC";
end if;
if pc = 17784 then
	inst <= x"002A0000";
end if;
if pc = 17788 then
	inst <= x"03DC0030";
end if;
if pc = 17792 then
	inst <= x"037E000C";
end if;
if pc = 17796 then
	inst <= x"C57DFFFC";
end if;
if pc = 17800 then
	inst <= x"8200400C";
end if;
if pc = 17804 then
	inst <= x"07DC0030";
end if;
if pc = 17808 then
	inst <= x"C05C0024";
end if;
if pc = 17812 then
	inst <= x"22640220";
end if;
if pc = 17816 then
	inst <= x"C09C0020";
end if;
if pc = 17820 then
	inst <= x"D4286000";
end if;
if pc = 17824 then
	inst <= x"820045D8";
end if;
if pc = 17828 then
	inst <= x"C49C0020";
end if;
if pc = 17832 then
	inst <= x"C43C0024";
end if;
if pc = 17836 then
	inst <= x"C17DFFFC";
end if;
if pc = 17840 then
	inst <= x"002A0000";
end if;
if pc = 17844 then
	inst <= x"03DC0030";
end if;
if pc = 17848 then
	inst <= x"037E000C";
end if;
if pc = 17852 then
	inst <= x"C57DFFFC";
end if;
if pc = 17856 then
	inst <= x"82003E98";
end if;
if pc = 17860 then
	inst <= x"07DC0030";
end if;
if pc = 17864 then
	inst <= x"C05C0024";
end if;
if pc = 17868 then
	inst <= x"22640220";
end if;
if pc = 17872 then
	inst <= x"C09C0020";
end if;
if pc = 17876 then
	inst <= x"D4286000";
end if;
if pc = 17880 then
	inst <= x"82004610";
end if;
if pc = 17884 then
	inst <= x"C49C0020";
end if;
if pc = 17888 then
	inst <= x"C43C0024";
end if;
if pc = 17892 then
	inst <= x"C17DFFFC";
end if;
if pc = 17896 then
	inst <= x"002A0000";
end if;
if pc = 17900 then
	inst <= x"03DC0030";
end if;
if pc = 17904 then
	inst <= x"037E000C";
end if;
if pc = 17908 then
	inst <= x"C57DFFFC";
end if;
if pc = 17912 then
	inst <= x"82003CC4";
end if;
if pc = 17916 then
	inst <= x"07DC0030";
end if;
if pc = 17920 then
	inst <= x"C05C0024";
end if;
if pc = 17924 then
	inst <= x"22640220";
end if;
if pc = 17928 then
	inst <= x"C09C0020";
end if;
if pc = 17932 then
	inst <= x"D4286000";
end if;
if pc = 17936 then
	inst <= x"06440001";
end if;
if pc = 17940 then
	inst <= x"C03C0000";
end if;
if pc = 17944 then
	inst <= x"820042A4";
end if;
if pc = 17948 then
	inst <= x"C1FDFFFC";
end if;
if pc = 17952 then
	inst <= x"C1FDFFFC";
end if;
if pc = 17956 then
	inst <= x"C1FDFFFC";
end if;
if pc = 17960 then
	inst <= x"C1FDFFFC";
end if;
if pc = 17964 then
	inst <= x"8640477C";
end if;
if pc = 17968 then
	inst <= x"026000C8";
end if;
if pc = 17972 then
	inst <= x"22840220";
end if;
if pc = 17976 then
	inst <= x"D0668000";
end if;
if pc = 17980 then
	inst <= x"C0860028";
end if;
if pc = 17984 then
	inst <= x"C0A60004";
end if;
if pc = 17988 then
	inst <= x"C8220000";
end if;
if pc = 17992 then
	inst <= x"C0C60014";
end if;
if pc = 17996 then
	inst <= x"C84C0000";
end if;
if pc = 18000 then
	inst <= x"44224000";
end if;
if pc = 18004 then
	inst <= x"CC280000";
end if;
if pc = 18008 then
	inst <= x"C8220004";
end if;
if pc = 18012 then
	inst <= x"C0C60014";
end if;
if pc = 18016 then
	inst <= x"C84C0004";
end if;
if pc = 18020 then
	inst <= x"44224000";
end if;
if pc = 18024 then
	inst <= x"CC280004";
end if;
if pc = 18028 then
	inst <= x"C8220008";
end if;
if pc = 18032 then
	inst <= x"C0C60014";
end if;
if pc = 18036 then
	inst <= x"C84C0008";
end if;
if pc = 18040 then
	inst <= x"44224000";
end if;
if pc = 18044 then
	inst <= x"CC280008";
end if;
if pc = 18048 then
	inst <= x"02C00002";
end if;
if pc = 18052 then
	inst <= x"82AC4740";
end if;
if pc = 18056 then
	inst <= x"02C00002";
end if;
if pc = 18060 then
	inst <= x"86CA4694";
end if;
if pc = 18064 then
	inst <= x"8200473C";
end if;
if pc = 18068 then
	inst <= x"C8280000";
end if;
if pc = 18072 then
	inst <= x"C8480004";
end if;
if pc = 18076 then
	inst <= x"C8680008";
end if;
if pc = 18080 then
	inst <= x"48822000";
end if;
if pc = 18084 then
	inst <= x"C0C60010";
end if;
if pc = 18088 then
	inst <= x"C8AC0000";
end if;
if pc = 18092 then
	inst <= x"4888A000";
end if;
if pc = 18096 then
	inst <= x"48A44000";
end if;
if pc = 18100 then
	inst <= x"C0C60010";
end if;
if pc = 18104 then
	inst <= x"C8CC0004";
end if;
if pc = 18108 then
	inst <= x"48AAC000";
end if;
if pc = 18112 then
	inst <= x"4088A000";
end if;
if pc = 18116 then
	inst <= x"48A66000";
end if;
if pc = 18120 then
	inst <= x"C0C60010";
end if;
if pc = 18124 then
	inst <= x"C8CC0008";
end if;
if pc = 18128 then
	inst <= x"48AAC000";
end if;
if pc = 18132 then
	inst <= x"4088A000";
end if;
if pc = 18136 then
	inst <= x"C0C6000C";
end if;
if pc = 18140 then
	inst <= x"82C04720";
end if;
if pc = 18144 then
	inst <= x"48A46000";
end if;
if pc = 18148 then
	inst <= x"C0C60024";
end if;
if pc = 18152 then
	inst <= x"C8CC0000";
end if;
if pc = 18156 then
	inst <= x"48AAC000";
end if;
if pc = 18160 then
	inst <= x"4088A000";
end if;
if pc = 18164 then
	inst <= x"48662000";
end if;
if pc = 18168 then
	inst <= x"C0C60024";
end if;
if pc = 18172 then
	inst <= x"C8AC0004";
end if;
if pc = 18176 then
	inst <= x"4866A000";
end if;
if pc = 18180 then
	inst <= x"40686000";
end if;
if pc = 18184 then
	inst <= x"48224000";
end if;
if pc = 18188 then
	inst <= x"C0660024";
end if;
if pc = 18192 then
	inst <= x"C8460008";
end if;
if pc = 18196 then
	inst <= x"48224000";
end if;
if pc = 18200 then
	inst <= x"40262000";
end if;
if pc = 18204 then
	inst <= x"82004724";
end if;
if pc = 18208 then
	inst <= x"40208000";
end if;
if pc = 18212 then
	inst <= x"02600003";
end if;
if pc = 18216 then
	inst <= x"82A64730";
end if;
if pc = 18220 then
	inst <= x"82004738";
end if;
if pc = 18224 then
	inst <= x"C84000A8";
end if;
if pc = 18228 then
	inst <= x"44224000";
end if;
if pc = 18232 then
	inst <= x"CC28000C";
end if;
if pc = 18236 then
	inst <= x"82004774";
end if;
if pc = 18240 then
	inst <= x"C0660010";
end if;
if pc = 18244 then
	inst <= x"C8280000";
end if;
if pc = 18248 then
	inst <= x"C8480004";
end if;
if pc = 18252 then
	inst <= x"C8680008";
end if;
if pc = 18256 then
	inst <= x"C8860000";
end if;
if pc = 18260 then
	inst <= x"48282000";
end if;
if pc = 18264 then
	inst <= x"C8860004";
end if;
if pc = 18268 then
	inst <= x"48484000";
end if;
if pc = 18272 then
	inst <= x"40224000";
end if;
if pc = 18276 then
	inst <= x"C8460008";
end if;
if pc = 18280 then
	inst <= x"48446000";
end if;
if pc = 18284 then
	inst <= x"40224000";
end if;
if pc = 18288 then
	inst <= x"CC28000C";
end if;
if pc = 18292 then
	inst <= x"06440001";
end if;
if pc = 18296 then
	inst <= x"8200462C";
end if;
if pc = 18300 then
	inst <= x"C1FDFFFC";
end if;
if pc = 18304 then
	inst <= x"48822000";
end if;
if pc = 18308 then
	inst <= x"C0420010";
end if;
if pc = 18312 then
	inst <= x"C8A40000";
end if;
if pc = 18316 then
	inst <= x"4888A000";
end if;
if pc = 18320 then
	inst <= x"48A44000";
end if;
if pc = 18324 then
	inst <= x"C0420010";
end if;
if pc = 18328 then
	inst <= x"C8C40004";
end if;
if pc = 18332 then
	inst <= x"48AAC000";
end if;
if pc = 18336 then
	inst <= x"4088A000";
end if;
if pc = 18340 then
	inst <= x"48A66000";
end if;
if pc = 18344 then
	inst <= x"C0420010";
end if;
if pc = 18348 then
	inst <= x"C8C40008";
end if;
if pc = 18352 then
	inst <= x"48AAC000";
end if;
if pc = 18356 then
	inst <= x"4088A000";
end if;
if pc = 18360 then
	inst <= x"C042000C";
end if;
if pc = 18364 then
	inst <= x"82404800";
end if;
if pc = 18368 then
	inst <= x"48A46000";
end if;
if pc = 18372 then
	inst <= x"C0420024";
end if;
if pc = 18376 then
	inst <= x"C8C40000";
end if;
if pc = 18380 then
	inst <= x"48AAC000";
end if;
if pc = 18384 then
	inst <= x"4088A000";
end if;
if pc = 18388 then
	inst <= x"48662000";
end if;
if pc = 18392 then
	inst <= x"C0420024";
end if;
if pc = 18396 then
	inst <= x"C8A40004";
end if;
if pc = 18400 then
	inst <= x"4866A000";
end if;
if pc = 18404 then
	inst <= x"40686000";
end if;
if pc = 18408 then
	inst <= x"48224000";
end if;
if pc = 18412 then
	inst <= x"C0420024";
end if;
if pc = 18416 then
	inst <= x"C8440008";
end if;
if pc = 18420 then
	inst <= x"48224000";
end if;
if pc = 18424 then
	inst <= x"40262000";
end if;
if pc = 18428 then
	inst <= x"82004804";
end if;
if pc = 18432 then
	inst <= x"40208000";
end if;
if pc = 18436 then
	inst <= x"C0420004";
end if;
if pc = 18440 then
	inst <= x"02600003";
end if;
if pc = 18444 then
	inst <= x"82464814";
end if;
if pc = 18448 then
	inst <= x"8200481C";
end if;
if pc = 18452 then
	inst <= x"C84000A8";
end if;
if pc = 18456 then
	inst <= x"44224000";
end if;
if pc = 18460 then
	inst <= x"C0220018";
end if;
if pc = 18464 then
	inst <= x"8E20482C";
end if;
if pc = 18468 then
	inst <= x"02400000";
end if;
if pc = 18472 then
	inst <= x"82004830";
end if;
if pc = 18476 then
	inst <= x"02400001";
end if;
if pc = 18480 then
	inst <= x"82204848";
end if;
if pc = 18484 then
	inst <= x"8E204840";
end if;
if pc = 18488 then
	inst <= x"02200001";
end if;
if pc = 18492 then
	inst <= x"82004844";
end if;
if pc = 18496 then
	inst <= x"02200000";
end if;
if pc = 18500 then
	inst <= x"8200484C";
end if;
if pc = 18504 then
	inst <= x"00240000";
end if;
if pc = 18508 then
	inst <= x"82204858";
end if;
if pc = 18512 then
	inst <= x"02200000";
end if;
if pc = 18516 then
	inst <= x"C1FDFFFC";
end if;
if pc = 18520 then
	inst <= x"02200001";
end if;
if pc = 18524 then
	inst <= x"C1FDFFFC";
end if;
if pc = 18528 then
	inst <= x"C0420014";
end if;
if pc = 18532 then
	inst <= x"C8840000";
end if;
if pc = 18536 then
	inst <= x"44228000";
end if;
if pc = 18540 then
	inst <= x"C0420014";
end if;
if pc = 18544 then
	inst <= x"C8840004";
end if;
if pc = 18548 then
	inst <= x"44448000";
end if;
if pc = 18552 then
	inst <= x"C0420014";
end if;
if pc = 18556 then
	inst <= x"C8840008";
end if;
if pc = 18560 then
	inst <= x"44668000";
end if;
if pc = 18564 then
	inst <= x"C0420004";
end if;
if pc = 18568 then
	inst <= x"02600001";
end if;
if pc = 18572 then
	inst <= x"8246497C";
end if;
if pc = 18576 then
	inst <= x"02600002";
end if;
if pc = 18580 then
	inst <= x"82464914";
end if;
if pc = 18584 then
	inst <= x"C43C0000";
end if;
if pc = 18588 then
	inst <= x"C17DFFFC";
end if;
if pc = 18592 then
	inst <= x"03DC000C";
end if;
if pc = 18596 then
	inst <= x"037E000C";
end if;
if pc = 18600 then
	inst <= x"C57DFFFC";
end if;
if pc = 18604 then
	inst <= x"82003344";
end if;
if pc = 18608 then
	inst <= x"07DC000C";
end if;
if pc = 18612 then
	inst <= x"C03C0000";
end if;
if pc = 18616 then
	inst <= x"C0420004";
end if;
if pc = 18620 then
	inst <= x"02600003";
end if;
if pc = 18624 then
	inst <= x"824648C8";
end if;
if pc = 18628 then
	inst <= x"820048D0";
end if;
if pc = 18632 then
	inst <= x"C84000A8";
end if;
if pc = 18636 then
	inst <= x"44224000";
end if;
if pc = 18640 then
	inst <= x"C0220018";
end if;
if pc = 18644 then
	inst <= x"8E2048E0";
end if;
if pc = 18648 then
	inst <= x"02400000";
end if;
if pc = 18652 then
	inst <= x"820048E4";
end if;
if pc = 18656 then
	inst <= x"02400001";
end if;
if pc = 18660 then
	inst <= x"822048FC";
end if;
if pc = 18664 then
	inst <= x"8E2048F4";
end if;
if pc = 18668 then
	inst <= x"02200001";
end if;
if pc = 18672 then
	inst <= x"820048F8";
end if;
if pc = 18676 then
	inst <= x"02200000";
end if;
if pc = 18680 then
	inst <= x"82004900";
end if;
if pc = 18684 then
	inst <= x"00240000";
end if;
if pc = 18688 then
	inst <= x"8220490C";
end if;
if pc = 18692 then
	inst <= x"02200000";
end if;
if pc = 18696 then
	inst <= x"C1FDFFFC";
end if;
if pc = 18700 then
	inst <= x"02200001";
end if;
if pc = 18704 then
	inst <= x"C1FDFFFC";
end if;
if pc = 18708 then
	inst <= x"C0420010";
end if;
if pc = 18712 then
	inst <= x"C8840000";
end if;
if pc = 18716 then
	inst <= x"48282000";
end if;
if pc = 18720 then
	inst <= x"C8840004";
end if;
if pc = 18724 then
	inst <= x"48484000";
end if;
if pc = 18728 then
	inst <= x"40224000";
end if;
if pc = 18732 then
	inst <= x"C8440008";
end if;
if pc = 18736 then
	inst <= x"48446000";
end if;
if pc = 18740 then
	inst <= x"40224000";
end if;
if pc = 18744 then
	inst <= x"C0220018";
end if;
if pc = 18748 then
	inst <= x"8E204948";
end if;
if pc = 18752 then
	inst <= x"02400000";
end if;
if pc = 18756 then
	inst <= x"8200494C";
end if;
if pc = 18760 then
	inst <= x"02400001";
end if;
if pc = 18764 then
	inst <= x"82204964";
end if;
if pc = 18768 then
	inst <= x"8E20495C";
end if;
if pc = 18772 then
	inst <= x"02200001";
end if;
if pc = 18776 then
	inst <= x"82004960";
end if;
if pc = 18780 then
	inst <= x"02200000";
end if;
if pc = 18784 then
	inst <= x"82004968";
end if;
if pc = 18788 then
	inst <= x"00240000";
end if;
if pc = 18792 then
	inst <= x"82204974";
end if;
if pc = 18796 then
	inst <= x"02200000";
end if;
if pc = 18800 then
	inst <= x"C1FDFFFC";
end if;
if pc = 18804 then
	inst <= x"02200001";
end if;
if pc = 18808 then
	inst <= x"C1FDFFFC";
end if;
if pc = 18812 then
	inst <= x"8E204984";
end if;
if pc = 18816 then
	inst <= x"82004988";
end if;
if pc = 18820 then
	inst <= x"44202000";
end if;
if pc = 18824 then
	inst <= x"C0420010";
end if;
if pc = 18828 then
	inst <= x"C8840000";
end if;
if pc = 18832 then
	inst <= x"8E28499C";
end if;
if pc = 18836 then
	inst <= x"02400000";
end if;
if pc = 18840 then
	inst <= x"820049E8";
end if;
if pc = 18844 then
	inst <= x"8E4049A8";
end if;
if pc = 18848 then
	inst <= x"40204000";
end if;
if pc = 18852 then
	inst <= x"820049AC";
end if;
if pc = 18856 then
	inst <= x"44204000";
end if;
if pc = 18860 then
	inst <= x"C0420010";
end if;
if pc = 18864 then
	inst <= x"C8440004";
end if;
if pc = 18868 then
	inst <= x"8E2449C0";
end if;
if pc = 18872 then
	inst <= x"02400000";
end if;
if pc = 18876 then
	inst <= x"820049E8";
end if;
if pc = 18880 then
	inst <= x"8E6049CC";
end if;
if pc = 18884 then
	inst <= x"40206000";
end if;
if pc = 18888 then
	inst <= x"820049D0";
end if;
if pc = 18892 then
	inst <= x"44206000";
end if;
if pc = 18896 then
	inst <= x"C0420010";
end if;
if pc = 18900 then
	inst <= x"C8440008";
end if;
if pc = 18904 then
	inst <= x"8E2449E4";
end if;
if pc = 18908 then
	inst <= x"02400000";
end if;
if pc = 18912 then
	inst <= x"820049E8";
end if;
if pc = 18916 then
	inst <= x"02400001";
end if;
if pc = 18920 then
	inst <= x"824049F4";
end if;
if pc = 18924 then
	inst <= x"C0220018";
end if;
if pc = 18928 then
	inst <= x"C1FDFFFC";
end if;
if pc = 18932 then
	inst <= x"C0220018";
end if;
if pc = 18936 then
	inst <= x"82204A04";
end if;
if pc = 18940 then
	inst <= x"02200000";
end if;
if pc = 18944 then
	inst <= x"C1FDFFFC";
end if;
if pc = 18948 then
	inst <= x"02200001";
end if;
if pc = 18952 then
	inst <= x"C1FDFFFC";
end if;
if pc = 18956 then
	inst <= x"22620220";
end if;
if pc = 18960 then
	inst <= x"D0646000";
end if;
if pc = 18964 then
	inst <= x"0280FFFF";
end if;
if pc = 18968 then
	inst <= x"82684E38";
end if;
if pc = 18972 then
	inst <= x"028000C8";
end if;
if pc = 18976 then
	inst <= x"22660220";
end if;
if pc = 18980 then
	inst <= x"D0686000";
end if;
if pc = 18984 then
	inst <= x"C0A60014";
end if;
if pc = 18988 then
	inst <= x"C88A0000";
end if;
if pc = 18992 then
	inst <= x"44828000";
end if;
if pc = 18996 then
	inst <= x"C0A60014";
end if;
if pc = 19000 then
	inst <= x"C8AA0004";
end if;
if pc = 19004 then
	inst <= x"44A4A000";
end if;
if pc = 19008 then
	inst <= x"C0A60014";
end if;
if pc = 19012 then
	inst <= x"C8CA0008";
end if;
if pc = 19016 then
	inst <= x"44C6C000";
end if;
if pc = 19020 then
	inst <= x"C0A60004";
end if;
if pc = 19024 then
	inst <= x"02C00001";
end if;
if pc = 19028 then
	inst <= x"CC7C0000";
end if;
if pc = 19032 then
	inst <= x"CC5C0008";
end if;
if pc = 19036 then
	inst <= x"CC3C0010";
end if;
if pc = 19040 then
	inst <= x"C49C0018";
end if;
if pc = 19044 then
	inst <= x"C45C001C";
end if;
if pc = 19048 then
	inst <= x"C43C0020";
end if;
if pc = 19052 then
	inst <= x"82AC4B0C";
end if;
if pc = 19056 then
	inst <= x"02C00002";
end if;
if pc = 19060 then
	inst <= x"82AC4AA4";
end if;
if pc = 19064 then
	inst <= x"C17DFFFC";
end if;
if pc = 19068 then
	inst <= x"00260000";
end if;
if pc = 19072 then
	inst <= x"4060C000";
end if;
if pc = 19076 then
	inst <= x"4040A000";
end if;
if pc = 19080 then
	inst <= x"40208000";
end if;
if pc = 19084 then
	inst <= x"03DC002C";
end if;
if pc = 19088 then
	inst <= x"037E000C";
end if;
if pc = 19092 then
	inst <= x"C57DFFFC";
end if;
if pc = 19096 then
	inst <= x"82004780";
end if;
if pc = 19100 then
	inst <= x"07DC002C";
end if;
if pc = 19104 then
	inst <= x"82004B08";
end if;
if pc = 19108 then
	inst <= x"C0A60010";
end if;
if pc = 19112 then
	inst <= x"C8EA0000";
end if;
if pc = 19116 then
	inst <= x"488E8000";
end if;
if pc = 19120 then
	inst <= x"C8EA0004";
end if;
if pc = 19124 then
	inst <= x"48AEA000";
end if;
if pc = 19128 then
	inst <= x"4088A000";
end if;
if pc = 19132 then
	inst <= x"C8AA0008";
end if;
if pc = 19136 then
	inst <= x"48AAC000";
end if;
if pc = 19140 then
	inst <= x"4088A000";
end if;
if pc = 19144 then
	inst <= x"C0660018";
end if;
if pc = 19148 then
	inst <= x"8E804AD8";
end if;
if pc = 19152 then
	inst <= x"02A00000";
end if;
if pc = 19156 then
	inst <= x"82004ADC";
end if;
if pc = 19160 then
	inst <= x"02A00001";
end if;
if pc = 19164 then
	inst <= x"82604AF4";
end if;
if pc = 19168 then
	inst <= x"8E804AEC";
end if;
if pc = 19172 then
	inst <= x"02600001";
end if;
if pc = 19176 then
	inst <= x"82004AF0";
end if;
if pc = 19180 then
	inst <= x"02600000";
end if;
if pc = 19184 then
	inst <= x"82004AF8";
end if;
if pc = 19188 then
	inst <= x"006A0000";
end if;
if pc = 19192 then
	inst <= x"82604B04";
end if;
if pc = 19196 then
	inst <= x"02200000";
end if;
if pc = 19200 then
	inst <= x"82004B08";
end if;
if pc = 19204 then
	inst <= x"02200001";
end if;
if pc = 19208 then
	inst <= x"82004B9C";
end if;
if pc = 19212 then
	inst <= x"8E804B14";
end if;
if pc = 19216 then
	inst <= x"82004B18";
end if;
if pc = 19220 then
	inst <= x"44808000";
end if;
if pc = 19224 then
	inst <= x"C0A60010";
end if;
if pc = 19228 then
	inst <= x"C8EA0000";
end if;
if pc = 19232 then
	inst <= x"8E8E4B2C";
end if;
if pc = 19236 then
	inst <= x"02A00000";
end if;
if pc = 19240 then
	inst <= x"82004B78";
end if;
if pc = 19244 then
	inst <= x"8EA04B38";
end if;
if pc = 19248 then
	inst <= x"4080A000";
end if;
if pc = 19252 then
	inst <= x"82004B3C";
end if;
if pc = 19256 then
	inst <= x"4480A000";
end if;
if pc = 19260 then
	inst <= x"C0A60010";
end if;
if pc = 19264 then
	inst <= x"C8AA0004";
end if;
if pc = 19268 then
	inst <= x"8E8A4B50";
end if;
if pc = 19272 then
	inst <= x"02A00000";
end if;
if pc = 19276 then
	inst <= x"82004B78";
end if;
if pc = 19280 then
	inst <= x"8EC04B5C";
end if;
if pc = 19284 then
	inst <= x"4080C000";
end if;
if pc = 19288 then
	inst <= x"82004B60";
end if;
if pc = 19292 then
	inst <= x"4480C000";
end if;
if pc = 19296 then
	inst <= x"C0A60010";
end if;
if pc = 19300 then
	inst <= x"C8AA0008";
end if;
if pc = 19304 then
	inst <= x"8E8A4B74";
end if;
if pc = 19308 then
	inst <= x"02A00000";
end if;
if pc = 19312 then
	inst <= x"82004B78";
end if;
if pc = 19316 then
	inst <= x"02A00001";
end if;
if pc = 19320 then
	inst <= x"82A04B88";
end if;
if pc = 19324 then
	inst <= x"C0660018";
end if;
if pc = 19328 then
	inst <= x"00260000";
end if;
if pc = 19332 then
	inst <= x"82004B9C";
end if;
if pc = 19336 then
	inst <= x"C0660018";
end if;
if pc = 19340 then
	inst <= x"82604B98";
end if;
if pc = 19344 then
	inst <= x"02200000";
end if;
if pc = 19348 then
	inst <= x"82004B9C";
end if;
if pc = 19352 then
	inst <= x"02200001";
end if;
if pc = 19356 then
	inst <= x"82204BA8";
end if;
if pc = 19360 then
	inst <= x"02200000";
end if;
if pc = 19364 then
	inst <= x"C1FDFFFC";
end if;
if pc = 19368 then
	inst <= x"C03C0020";
end if;
if pc = 19372 then
	inst <= x"02220001";
end if;
if pc = 19376 then
	inst <= x"22420220";
end if;
if pc = 19380 then
	inst <= x"C07C001C";
end if;
if pc = 19384 then
	inst <= x"D0464000";
end if;
if pc = 19388 then
	inst <= x"0280FFFF";
end if;
if pc = 19392 then
	inst <= x"82484E30";
end if;
if pc = 19396 then
	inst <= x"22440220";
end if;
if pc = 19400 then
	inst <= x"C09C0018";
end if;
if pc = 19404 then
	inst <= x"D0484000";
end if;
if pc = 19408 then
	inst <= x"C83C0010";
end if;
if pc = 19412 then
	inst <= x"C85C0008";
end if;
if pc = 19416 then
	inst <= x"C87C0000";
end if;
if pc = 19420 then
	inst <= x"C43C0024";
end if;
if pc = 19424 then
	inst <= x"C17DFFFC";
end if;
if pc = 19428 then
	inst <= x"00240000";
end if;
if pc = 19432 then
	inst <= x"03DC0030";
end if;
if pc = 19436 then
	inst <= x"037E000C";
end if;
if pc = 19440 then
	inst <= x"C57DFFFC";
end if;
if pc = 19444 then
	inst <= x"82004860";
end if;
if pc = 19448 then
	inst <= x"07DC0030";
end if;
if pc = 19452 then
	inst <= x"82204C08";
end if;
if pc = 19456 then
	inst <= x"02200000";
end if;
if pc = 19460 then
	inst <= x"C1FDFFFC";
end if;
if pc = 19464 then
	inst <= x"C03C0024";
end if;
if pc = 19468 then
	inst <= x"02220001";
end if;
if pc = 19472 then
	inst <= x"22420220";
end if;
if pc = 19476 then
	inst <= x"C07C001C";
end if;
if pc = 19480 then
	inst <= x"D0464000";
end if;
if pc = 19484 then
	inst <= x"0280FFFF";
end if;
if pc = 19488 then
	inst <= x"82484E28";
end if;
if pc = 19492 then
	inst <= x"22440220";
end if;
if pc = 19496 then
	inst <= x"C09C0018";
end if;
if pc = 19500 then
	inst <= x"D0484000";
end if;
if pc = 19504 then
	inst <= x"C0A40014";
end if;
if pc = 19508 then
	inst <= x"C82A0000";
end if;
if pc = 19512 then
	inst <= x"C85C0010";
end if;
if pc = 19516 then
	inst <= x"44242000";
end if;
if pc = 19520 then
	inst <= x"C0A40014";
end if;
if pc = 19524 then
	inst <= x"C86A0004";
end if;
if pc = 19528 then
	inst <= x"C89C0008";
end if;
if pc = 19532 then
	inst <= x"44686000";
end if;
if pc = 19536 then
	inst <= x"C0A40014";
end if;
if pc = 19540 then
	inst <= x"C8AA0008";
end if;
if pc = 19544 then
	inst <= x"C8DC0000";
end if;
if pc = 19548 then
	inst <= x"44ACA000";
end if;
if pc = 19552 then
	inst <= x"C0A40004";
end if;
if pc = 19556 then
	inst <= x"02C00001";
end if;
if pc = 19560 then
	inst <= x"C43C0028";
end if;
if pc = 19564 then
	inst <= x"82AC4D08";
end if;
if pc = 19568 then
	inst <= x"02C00002";
end if;
if pc = 19572 then
	inst <= x"82AC4CA0";
end if;
if pc = 19576 then
	inst <= x"C17DFFFC";
end if;
if pc = 19580 then
	inst <= x"00240000";
end if;
if pc = 19584 then
	inst <= x"40406000";
end if;
if pc = 19588 then
	inst <= x"4060A000";
end if;
if pc = 19592 then
	inst <= x"03DC0034";
end if;
if pc = 19596 then
	inst <= x"037E000C";
end if;
if pc = 19600 then
	inst <= x"C57DFFFC";
end if;
if pc = 19604 then
	inst <= x"82004780";
end if;
if pc = 19608 then
	inst <= x"07DC0034";
end if;
if pc = 19612 then
	inst <= x"82004D04";
end if;
if pc = 19616 then
	inst <= x"C0A40010";
end if;
if pc = 19620 then
	inst <= x"C8EA0000";
end if;
if pc = 19624 then
	inst <= x"482E2000";
end if;
if pc = 19628 then
	inst <= x"C8EA0004";
end if;
if pc = 19632 then
	inst <= x"486E6000";
end if;
if pc = 19636 then
	inst <= x"40226000";
end if;
if pc = 19640 then
	inst <= x"C86A0008";
end if;
if pc = 19644 then
	inst <= x"4866A000";
end if;
if pc = 19648 then
	inst <= x"40226000";
end if;
if pc = 19652 then
	inst <= x"C0440018";
end if;
if pc = 19656 then
	inst <= x"8E204CD4";
end if;
if pc = 19660 then
	inst <= x"02A00000";
end if;
if pc = 19664 then
	inst <= x"82004CD8";
end if;
if pc = 19668 then
	inst <= x"02A00001";
end if;
if pc = 19672 then
	inst <= x"82404CF0";
end if;
if pc = 19676 then
	inst <= x"8E204CE8";
end if;
if pc = 19680 then
	inst <= x"02400001";
end if;
if pc = 19684 then
	inst <= x"82004CEC";
end if;
if pc = 19688 then
	inst <= x"02400000";
end if;
if pc = 19692 then
	inst <= x"82004CF4";
end if;
if pc = 19696 then
	inst <= x"004A0000";
end if;
if pc = 19700 then
	inst <= x"82404D00";
end if;
if pc = 19704 then
	inst <= x"02200000";
end if;
if pc = 19708 then
	inst <= x"82004D04";
end if;
if pc = 19712 then
	inst <= x"02200001";
end if;
if pc = 19716 then
	inst <= x"82004D98";
end if;
if pc = 19720 then
	inst <= x"8E204D10";
end if;
if pc = 19724 then
	inst <= x"82004D14";
end if;
if pc = 19728 then
	inst <= x"44202000";
end if;
if pc = 19732 then
	inst <= x"C0A40010";
end if;
if pc = 19736 then
	inst <= x"C8EA0000";
end if;
if pc = 19740 then
	inst <= x"8E2E4D28";
end if;
if pc = 19744 then
	inst <= x"02A00000";
end if;
if pc = 19748 then
	inst <= x"82004D74";
end if;
if pc = 19752 then
	inst <= x"8E604D34";
end if;
if pc = 19756 then
	inst <= x"40206000";
end if;
if pc = 19760 then
	inst <= x"82004D38";
end if;
if pc = 19764 then
	inst <= x"44206000";
end if;
if pc = 19768 then
	inst <= x"C0A40010";
end if;
if pc = 19772 then
	inst <= x"C86A0004";
end if;
if pc = 19776 then
	inst <= x"8E264D4C";
end if;
if pc = 19780 then
	inst <= x"02A00000";
end if;
if pc = 19784 then
	inst <= x"82004D74";
end if;
if pc = 19788 then
	inst <= x"8EA04D58";
end if;
if pc = 19792 then
	inst <= x"4020A000";
end if;
if pc = 19796 then
	inst <= x"82004D5C";
end if;
if pc = 19800 then
	inst <= x"4420A000";
end if;
if pc = 19804 then
	inst <= x"C0A40010";
end if;
if pc = 19808 then
	inst <= x"C86A0008";
end if;
if pc = 19812 then
	inst <= x"8E264D70";
end if;
if pc = 19816 then
	inst <= x"02A00000";
end if;
if pc = 19820 then
	inst <= x"82004D74";
end if;
if pc = 19824 then
	inst <= x"02A00001";
end if;
if pc = 19828 then
	inst <= x"82A04D84";
end if;
if pc = 19832 then
	inst <= x"C0440018";
end if;
if pc = 19836 then
	inst <= x"00240000";
end if;
if pc = 19840 then
	inst <= x"82004D98";
end if;
if pc = 19844 then
	inst <= x"C0440018";
end if;
if pc = 19848 then
	inst <= x"82404D94";
end if;
if pc = 19852 then
	inst <= x"02200000";
end if;
if pc = 19856 then
	inst <= x"82004D98";
end if;
if pc = 19860 then
	inst <= x"02200001";
end if;
if pc = 19864 then
	inst <= x"82204DA4";
end if;
if pc = 19868 then
	inst <= x"02200000";
end if;
if pc = 19872 then
	inst <= x"C1FDFFFC";
end if;
if pc = 19876 then
	inst <= x"C03C0028";
end if;
if pc = 19880 then
	inst <= x"02220001";
end if;
if pc = 19884 then
	inst <= x"22420220";
end if;
if pc = 19888 then
	inst <= x"C07C001C";
end if;
if pc = 19892 then
	inst <= x"D0464000";
end if;
if pc = 19896 then
	inst <= x"0280FFFF";
end if;
if pc = 19900 then
	inst <= x"82484E20";
end if;
if pc = 19904 then
	inst <= x"22440220";
end if;
if pc = 19908 then
	inst <= x"C09C0018";
end if;
if pc = 19912 then
	inst <= x"D0484000";
end if;
if pc = 19916 then
	inst <= x"C83C0010";
end if;
if pc = 19920 then
	inst <= x"C85C0008";
end if;
if pc = 19924 then
	inst <= x"C87C0000";
end if;
if pc = 19928 then
	inst <= x"C43C002C";
end if;
if pc = 19932 then
	inst <= x"C17DFFFC";
end if;
if pc = 19936 then
	inst <= x"00240000";
end if;
if pc = 19940 then
	inst <= x"03DC0038";
end if;
if pc = 19944 then
	inst <= x"037E000C";
end if;
if pc = 19948 then
	inst <= x"C57DFFFC";
end if;
if pc = 19952 then
	inst <= x"82004860";
end if;
if pc = 19956 then
	inst <= x"07DC0038";
end if;
if pc = 19960 then
	inst <= x"82204E04";
end if;
if pc = 19964 then
	inst <= x"02200000";
end if;
if pc = 19968 then
	inst <= x"C1FDFFFC";
end if;
if pc = 19972 then
	inst <= x"C03C002C";
end if;
if pc = 19976 then
	inst <= x"02220001";
end if;
if pc = 19980 then
	inst <= x"C83C0010";
end if;
if pc = 19984 then
	inst <= x"C85C0008";
end if;
if pc = 19988 then
	inst <= x"C87C0000";
end if;
if pc = 19992 then
	inst <= x"C05C001C";
end if;
if pc = 19996 then
	inst <= x"82004A0C";
end if;
if pc = 20000 then
	inst <= x"02200001";
end if;
if pc = 20004 then
	inst <= x"C1FDFFFC";
end if;
if pc = 20008 then
	inst <= x"02200001";
end if;
if pc = 20012 then
	inst <= x"C1FDFFFC";
end if;
if pc = 20016 then
	inst <= x"02200001";
end if;
if pc = 20020 then
	inst <= x"C1FDFFFC";
end if;
if pc = 20024 then
	inst <= x"02200001";
end if;
if pc = 20028 then
	inst <= x"C1FDFFFC";
end if;
if pc = 20032 then
	inst <= x"22620220";
end if;
if pc = 20036 then
	inst <= x"D0646000";
end if;
if pc = 20040 then
	inst <= x"0280FFFF";
end if;
if pc = 20044 then
	inst <= x"8268527C";
end if;
if pc = 20048 then
	inst <= x"02800368";
end if;
if pc = 20052 then
	inst <= x"02A002B8";
end if;
if pc = 20056 then
	inst <= x"02C000C8";
end if;
if pc = 20060 then
	inst <= x"22E60220";
end if;
if pc = 20064 then
	inst <= x"D0ECE000";
end if;
if pc = 20068 then
	inst <= x"C82A0000";
end if;
if pc = 20072 then
	inst <= x"C10E0014";
end if;
if pc = 20076 then
	inst <= x"C8500000";
end if;
if pc = 20080 then
	inst <= x"44224000";
end if;
if pc = 20084 then
	inst <= x"C84A0004";
end if;
if pc = 20088 then
	inst <= x"C10E0014";
end if;
if pc = 20092 then
	inst <= x"C8700004";
end if;
if pc = 20096 then
	inst <= x"44446000";
end if;
if pc = 20100 then
	inst <= x"C86A0008";
end if;
if pc = 20104 then
	inst <= x"C10E0014";
end if;
if pc = 20108 then
	inst <= x"C8900008";
end if;
if pc = 20112 then
	inst <= x"44668000";
end if;
if pc = 20116 then
	inst <= x"C1080004";
end if;
if pc = 20120 then
	inst <= x"23260220";
end if;
if pc = 20124 then
	inst <= x"D1112000";
end if;
if pc = 20128 then
	inst <= x"C12E0004";
end if;
if pc = 20132 then
	inst <= x"03400001";
end if;
if pc = 20136 then
	inst <= x"C4BC0000";
end if;
if pc = 20140 then
	inst <= x"C45C0004";
end if;
if pc = 20144 then
	inst <= x"C43C0008";
end if;
if pc = 20148 then
	inst <= x"C4DC000C";
end if;
if pc = 20152 then
	inst <= x"C47C0010";
end if;
if pc = 20156 then
	inst <= x"83344F2C";
end if;
if pc = 20160 then
	inst <= x"02800002";
end if;
if pc = 20164 then
	inst <= x"83284EEC";
end if;
if pc = 20168 then
	inst <= x"C17DFFFC";
end if;
if pc = 20172 then
	inst <= x"00500000";
end if;
if pc = 20176 then
	inst <= x"002E0000";
end if;
if pc = 20180 then
	inst <= x"03DC001C";
end if;
if pc = 20184 then
	inst <= x"037E000C";
end if;
if pc = 20188 then
	inst <= x"C57DFFFC";
end if;
if pc = 20192 then
	inst <= x"82003A54";
end if;
if pc = 20196 then
	inst <= x"07DC001C";
end if;
if pc = 20200 then
	inst <= x"82004F28";
end if;
if pc = 20204 then
	inst <= x"C8900000";
end if;
if pc = 20208 then
	inst <= x"8E804EFC";
end if;
if pc = 20212 then
	inst <= x"02200000";
end if;
if pc = 20216 then
	inst <= x"82004F28";
end if;
if pc = 20220 then
	inst <= x"028002AC";
end if;
if pc = 20224 then
	inst <= x"C8900004";
end if;
if pc = 20228 then
	inst <= x"48282000";
end if;
if pc = 20232 then
	inst <= x"C8900008";
end if;
if pc = 20236 then
	inst <= x"48484000";
end if;
if pc = 20240 then
	inst <= x"40224000";
end if;
if pc = 20244 then
	inst <= x"C850000C";
end if;
if pc = 20248 then
	inst <= x"48446000";
end if;
if pc = 20252 then
	inst <= x"40224000";
end if;
if pc = 20256 then
	inst <= x"CC280000";
end if;
if pc = 20260 then
	inst <= x"02200001";
end if;
if pc = 20264 then
	inst <= x"82004F54";
end if;
if pc = 20268 then
	inst <= x"C0880000";
end if;
if pc = 20272 then
	inst <= x"C17DFFFC";
end if;
if pc = 20276 then
	inst <= x"00700000";
end if;
if pc = 20280 then
	inst <= x"00480000";
end if;
if pc = 20284 then
	inst <= x"002E0000";
end if;
if pc = 20288 then
	inst <= x"03DC001C";
end if;
if pc = 20292 then
	inst <= x"037E000C";
end if;
if pc = 20296 then
	inst <= x"C57DFFFC";
end if;
if pc = 20300 then
	inst <= x"8200389C";
end if;
if pc = 20304 then
	inst <= x"07DC001C";
end if;
if pc = 20308 then
	inst <= x"024002AC";
end if;
if pc = 20312 then
	inst <= x"C8240000";
end if;
if pc = 20316 then
	inst <= x"82204F78";
end if;
if pc = 20320 then
	inst <= x"C8400078";
end if;
if pc = 20324 then
	inst <= x"8E244F70";
end if;
if pc = 20328 then
	inst <= x"02200000";
end if;
if pc = 20332 then
	inst <= x"82004F74";
end if;
if pc = 20336 then
	inst <= x"02200001";
end if;
if pc = 20340 then
	inst <= x"82004F7C";
end if;
if pc = 20344 then
	inst <= x"02200000";
end if;
if pc = 20348 then
	inst <= x"8220524C";
end if;
if pc = 20352 then
	inst <= x"C8400074";
end if;
if pc = 20356 then
	inst <= x"40224000";
end if;
if pc = 20360 then
	inst <= x"022001D0";
end if;
if pc = 20364 then
	inst <= x"C8420000";
end if;
if pc = 20368 then
	inst <= x"48442000";
end if;
if pc = 20372 then
	inst <= x"C05C0000";
end if;
if pc = 20376 then
	inst <= x"C8640000";
end if;
if pc = 20380 then
	inst <= x"40446000";
end if;
if pc = 20384 then
	inst <= x"C8620004";
end if;
if pc = 20388 then
	inst <= x"48662000";
end if;
if pc = 20392 then
	inst <= x"C8840004";
end if;
if pc = 20396 then
	inst <= x"40668000";
end if;
if pc = 20400 then
	inst <= x"C8820008";
end if;
if pc = 20404 then
	inst <= x"48282000";
end if;
if pc = 20408 then
	inst <= x"C8840008";
end if;
if pc = 20412 then
	inst <= x"40228000";
end if;
if pc = 20416 then
	inst <= x"C05C0004";
end if;
if pc = 20420 then
	inst <= x"C0240000";
end if;
if pc = 20424 then
	inst <= x"0260FFFF";
end if;
if pc = 20428 then
	inst <= x"8226522C";
end if;
if pc = 20432 then
	inst <= x"22220220";
end if;
if pc = 20436 then
	inst <= x"C07C000C";
end if;
if pc = 20440 then
	inst <= x"D0262000";
end if;
if pc = 20444 then
	inst <= x"CC3C0018";
end if;
if pc = 20448 then
	inst <= x"CC7C0020";
end if;
if pc = 20452 then
	inst <= x"CC5C0028";
end if;
if pc = 20456 then
	inst <= x"C17DFFFC";
end if;
if pc = 20460 then
	inst <= x"41E06000";
end if;
if pc = 20464 then
	inst <= x"40602000";
end if;
if pc = 20468 then
	inst <= x"40204000";
end if;
if pc = 20472 then
	inst <= x"4041E000";
end if;
if pc = 20476 then
	inst <= x"03DC0038";
end if;
if pc = 20480 then
	inst <= x"037E000C";
end if;
if pc = 20484 then
	inst <= x"C57DFFFC";
end if;
if pc = 20488 then
	inst <= x"82004860";
end if;
if pc = 20492 then
	inst <= x"07DC0038";
end if;
if pc = 20496 then
	inst <= x"8220501C";
end if;
if pc = 20500 then
	inst <= x"02200000";
end if;
if pc = 20504 then
	inst <= x"82005228";
end if;
if pc = 20508 then
	inst <= x"C05C0004";
end if;
if pc = 20512 then
	inst <= x"C0240004";
end if;
if pc = 20516 then
	inst <= x"0260FFFF";
end if;
if pc = 20520 then
	inst <= x"82265224";
end if;
if pc = 20524 then
	inst <= x"22220220";
end if;
if pc = 20528 then
	inst <= x"C07C000C";
end if;
if pc = 20532 then
	inst <= x"D0262000";
end if;
if pc = 20536 then
	inst <= x"C0820014";
end if;
if pc = 20540 then
	inst <= x"C8280000";
end if;
if pc = 20544 then
	inst <= x"C85C0028";
end if;
if pc = 20548 then
	inst <= x"44242000";
end if;
if pc = 20552 then
	inst <= x"C0820014";
end if;
if pc = 20556 then
	inst <= x"C8680004";
end if;
if pc = 20560 then
	inst <= x"C89C0020";
end if;
if pc = 20564 then
	inst <= x"44686000";
end if;
if pc = 20568 then
	inst <= x"C0820014";
end if;
if pc = 20572 then
	inst <= x"C8A80008";
end if;
if pc = 20576 then
	inst <= x"C8DC0018";
end if;
if pc = 20580 then
	inst <= x"44ACA000";
end if;
if pc = 20584 then
	inst <= x"C0820004";
end if;
if pc = 20588 then
	inst <= x"02A00001";
end if;
if pc = 20592 then
	inst <= x"828A5108";
end if;
if pc = 20596 then
	inst <= x"02A00002";
end if;
if pc = 20600 then
	inst <= x"828A50A0";
end if;
if pc = 20604 then
	inst <= x"C17DFFFC";
end if;
if pc = 20608 then
	inst <= x"40406000";
end if;
if pc = 20612 then
	inst <= x"4060A000";
end if;
if pc = 20616 then
	inst <= x"03DC0038";
end if;
if pc = 20620 then
	inst <= x"037E000C";
end if;
if pc = 20624 then
	inst <= x"C57DFFFC";
end if;
if pc = 20628 then
	inst <= x"82004780";
end if;
if pc = 20632 then
	inst <= x"07DC0038";
end if;
if pc = 20636 then
	inst <= x"82005104";
end if;
if pc = 20640 then
	inst <= x"C0820010";
end if;
if pc = 20644 then
	inst <= x"C8E80000";
end if;
if pc = 20648 then
	inst <= x"482E2000";
end if;
if pc = 20652 then
	inst <= x"C8E80004";
end if;
if pc = 20656 then
	inst <= x"486E6000";
end if;
if pc = 20660 then
	inst <= x"40226000";
end if;
if pc = 20664 then
	inst <= x"C8680008";
end if;
if pc = 20668 then
	inst <= x"4866A000";
end if;
if pc = 20672 then
	inst <= x"40226000";
end if;
if pc = 20676 then
	inst <= x"C0220018";
end if;
if pc = 20680 then
	inst <= x"8E2050D4";
end if;
if pc = 20684 then
	inst <= x"02800000";
end if;
if pc = 20688 then
	inst <= x"820050D8";
end if;
if pc = 20692 then
	inst <= x"02800001";
end if;
if pc = 20696 then
	inst <= x"822050F0";
end if;
if pc = 20700 then
	inst <= x"8E2050E8";
end if;
if pc = 20704 then
	inst <= x"02200001";
end if;
if pc = 20708 then
	inst <= x"820050EC";
end if;
if pc = 20712 then
	inst <= x"02200000";
end if;
if pc = 20716 then
	inst <= x"820050F4";
end if;
if pc = 20720 then
	inst <= x"00280000";
end if;
if pc = 20724 then
	inst <= x"82205100";
end if;
if pc = 20728 then
	inst <= x"02200000";
end if;
if pc = 20732 then
	inst <= x"82005104";
end if;
if pc = 20736 then
	inst <= x"02200001";
end if;
if pc = 20740 then
	inst <= x"82005194";
end if;
if pc = 20744 then
	inst <= x"8E205110";
end if;
if pc = 20748 then
	inst <= x"82005114";
end if;
if pc = 20752 then
	inst <= x"44202000";
end if;
if pc = 20756 then
	inst <= x"C0820010";
end if;
if pc = 20760 then
	inst <= x"C8E80000";
end if;
if pc = 20764 then
	inst <= x"8E2E5128";
end if;
if pc = 20768 then
	inst <= x"02800000";
end if;
if pc = 20772 then
	inst <= x"82005174";
end if;
if pc = 20776 then
	inst <= x"8E605134";
end if;
if pc = 20780 then
	inst <= x"40206000";
end if;
if pc = 20784 then
	inst <= x"82005138";
end if;
if pc = 20788 then
	inst <= x"44206000";
end if;
if pc = 20792 then
	inst <= x"C0820010";
end if;
if pc = 20796 then
	inst <= x"C8680004";
end if;
if pc = 20800 then
	inst <= x"8E26514C";
end if;
if pc = 20804 then
	inst <= x"02800000";
end if;
if pc = 20808 then
	inst <= x"82005174";
end if;
if pc = 20812 then
	inst <= x"8EA05158";
end if;
if pc = 20816 then
	inst <= x"4020A000";
end if;
if pc = 20820 then
	inst <= x"8200515C";
end if;
if pc = 20824 then
	inst <= x"4420A000";
end if;
if pc = 20828 then
	inst <= x"C0820010";
end if;
if pc = 20832 then
	inst <= x"C8680008";
end if;
if pc = 20836 then
	inst <= x"8E265170";
end if;
if pc = 20840 then
	inst <= x"02800000";
end if;
if pc = 20844 then
	inst <= x"82005174";
end if;
if pc = 20848 then
	inst <= x"02800001";
end if;
if pc = 20852 then
	inst <= x"82805180";
end if;
if pc = 20856 then
	inst <= x"C0220018";
end if;
if pc = 20860 then
	inst <= x"82005194";
end if;
if pc = 20864 then
	inst <= x"C0220018";
end if;
if pc = 20868 then
	inst <= x"82205190";
end if;
if pc = 20872 then
	inst <= x"02200000";
end if;
if pc = 20876 then
	inst <= x"82005194";
end if;
if pc = 20880 then
	inst <= x"02200001";
end if;
if pc = 20884 then
	inst <= x"822051A0";
end if;
if pc = 20888 then
	inst <= x"02200000";
end if;
if pc = 20892 then
	inst <= x"82005220";
end if;
if pc = 20896 then
	inst <= x"C05C0004";
end if;
if pc = 20900 then
	inst <= x"C0240008";
end if;
if pc = 20904 then
	inst <= x"0260FFFF";
end if;
if pc = 20908 then
	inst <= x"8226521C";
end if;
if pc = 20912 then
	inst <= x"22220220";
end if;
if pc = 20916 then
	inst <= x"C07C000C";
end if;
if pc = 20920 then
	inst <= x"D0262000";
end if;
if pc = 20924 then
	inst <= x"C83C0028";
end if;
if pc = 20928 then
	inst <= x"C85C0020";
end if;
if pc = 20932 then
	inst <= x"C87C0018";
end if;
if pc = 20936 then
	inst <= x"C17DFFFC";
end if;
if pc = 20940 then
	inst <= x"03DC0038";
end if;
if pc = 20944 then
	inst <= x"037E000C";
end if;
if pc = 20948 then
	inst <= x"C57DFFFC";
end if;
if pc = 20952 then
	inst <= x"82004860";
end if;
if pc = 20956 then
	inst <= x"07DC0038";
end if;
if pc = 20960 then
	inst <= x"822051EC";
end if;
if pc = 20964 then
	inst <= x"02200000";
end if;
if pc = 20968 then
	inst <= x"82005218";
end if;
if pc = 20972 then
	inst <= x"02200003";
end if;
if pc = 20976 then
	inst <= x"C83C0028";
end if;
if pc = 20980 then
	inst <= x"C85C0020";
end if;
if pc = 20984 then
	inst <= x"C87C0018";
end if;
if pc = 20988 then
	inst <= x"C05C0004";
end if;
if pc = 20992 then
	inst <= x"C17DFFFC";
end if;
if pc = 20996 then
	inst <= x"03DC0038";
end if;
if pc = 21000 then
	inst <= x"037E000C";
end if;
if pc = 21004 then
	inst <= x"C57DFFFC";
end if;
if pc = 21008 then
	inst <= x"82004A0C";
end if;
if pc = 21012 then
	inst <= x"07DC0038";
end if;
if pc = 21016 then
	inst <= x"82005220";
end if;
if pc = 21020 then
	inst <= x"02200001";
end if;
if pc = 21024 then
	inst <= x"82005228";
end if;
if pc = 21028 then
	inst <= x"02200001";
end if;
if pc = 21032 then
	inst <= x"82005230";
end if;
if pc = 21036 then
	inst <= x"02200001";
end if;
if pc = 21040 then
	inst <= x"8220523C";
end if;
if pc = 21044 then
	inst <= x"02200001";
end if;
if pc = 21048 then
	inst <= x"C1FDFFFC";
end if;
if pc = 21052 then
	inst <= x"C03C0008";
end if;
if pc = 21056 then
	inst <= x"02220001";
end if;
if pc = 21060 then
	inst <= x"C05C0004";
end if;
if pc = 21064 then
	inst <= x"82004E40";
end if;
if pc = 21068 then
	inst <= x"C03C0010";
end if;
if pc = 21072 then
	inst <= x"22220220";
end if;
if pc = 21076 then
	inst <= x"C05C000C";
end if;
if pc = 21080 then
	inst <= x"D0242000";
end if;
if pc = 21084 then
	inst <= x"C0220018";
end if;
if pc = 21088 then
	inst <= x"82205274";
end if;
if pc = 21092 then
	inst <= x"C03C0008";
end if;
if pc = 21096 then
	inst <= x"02220001";
end if;
if pc = 21100 then
	inst <= x"C05C0004";
end if;
if pc = 21104 then
	inst <= x"82004E40";
end if;
if pc = 21108 then
	inst <= x"02200000";
end if;
if pc = 21112 then
	inst <= x"C1FDFFFC";
end if;
if pc = 21116 then
	inst <= x"02200000";
end if;
if pc = 21120 then
	inst <= x"C1FDFFFC";
end if;
if pc = 21124 then
	inst <= x"22620220";
end if;
if pc = 21128 then
	inst <= x"D0646000";
end if;
if pc = 21132 then
	inst <= x"0280FFFF";
end if;
if pc = 21136 then
	inst <= x"8268540C";
end if;
if pc = 21140 then
	inst <= x"028001E0";
end if;
if pc = 21144 then
	inst <= x"22660220";
end if;
if pc = 21148 then
	inst <= x"D0686000";
end if;
if pc = 21152 then
	inst <= x"02A00000";
end if;
if pc = 21156 then
	inst <= x"C49C0000";
end if;
if pc = 21160 then
	inst <= x"C45C0004";
end if;
if pc = 21164 then
	inst <= x"C43C0008";
end if;
if pc = 21168 then
	inst <= x"C17DFFFC";
end if;
if pc = 21172 then
	inst <= x"00460000";
end if;
if pc = 21176 then
	inst <= x"002A0000";
end if;
if pc = 21180 then
	inst <= x"03DC0014";
end if;
if pc = 21184 then
	inst <= x"037E000C";
end if;
if pc = 21188 then
	inst <= x"C57DFFFC";
end if;
if pc = 21192 then
	inst <= x"82004E40";
end if;
if pc = 21196 then
	inst <= x"07DC0014";
end if;
if pc = 21200 then
	inst <= x"822052DC";
end if;
if pc = 21204 then
	inst <= x"02200001";
end if;
if pc = 21208 then
	inst <= x"C1FDFFFC";
end if;
if pc = 21212 then
	inst <= x"C03C0008";
end if;
if pc = 21216 then
	inst <= x"02220001";
end if;
if pc = 21220 then
	inst <= x"22420220";
end if;
if pc = 21224 then
	inst <= x"C07C0004";
end if;
if pc = 21228 then
	inst <= x"D0464000";
end if;
if pc = 21232 then
	inst <= x"0280FFFF";
end if;
if pc = 21236 then
	inst <= x"82485404";
end if;
if pc = 21240 then
	inst <= x"22440220";
end if;
if pc = 21244 then
	inst <= x"C09C0000";
end if;
if pc = 21248 then
	inst <= x"D0484000";
end if;
if pc = 21252 then
	inst <= x"02A00000";
end if;
if pc = 21256 then
	inst <= x"C43C000C";
end if;
if pc = 21260 then
	inst <= x"C17DFFFC";
end if;
if pc = 21264 then
	inst <= x"002A0000";
end if;
if pc = 21268 then
	inst <= x"03DC0018";
end if;
if pc = 21272 then
	inst <= x"037E000C";
end if;
if pc = 21276 then
	inst <= x"C57DFFFC";
end if;
if pc = 21280 then
	inst <= x"82004E40";
end if;
if pc = 21284 then
	inst <= x"07DC0018";
end if;
if pc = 21288 then
	inst <= x"82205334";
end if;
if pc = 21292 then
	inst <= x"02200001";
end if;
if pc = 21296 then
	inst <= x"C1FDFFFC";
end if;
if pc = 21300 then
	inst <= x"C03C000C";
end if;
if pc = 21304 then
	inst <= x"02220001";
end if;
if pc = 21308 then
	inst <= x"22420220";
end if;
if pc = 21312 then
	inst <= x"C07C0004";
end if;
if pc = 21316 then
	inst <= x"D0464000";
end if;
if pc = 21320 then
	inst <= x"0280FFFF";
end if;
if pc = 21324 then
	inst <= x"824853FC";
end if;
if pc = 21328 then
	inst <= x"22440220";
end if;
if pc = 21332 then
	inst <= x"C09C0000";
end if;
if pc = 21336 then
	inst <= x"D0484000";
end if;
if pc = 21340 then
	inst <= x"02A00000";
end if;
if pc = 21344 then
	inst <= x"C43C0010";
end if;
if pc = 21348 then
	inst <= x"C17DFFFC";
end if;
if pc = 21352 then
	inst <= x"002A0000";
end if;
if pc = 21356 then
	inst <= x"03DC001C";
end if;
if pc = 21360 then
	inst <= x"037E000C";
end if;
if pc = 21364 then
	inst <= x"C57DFFFC";
end if;
if pc = 21368 then
	inst <= x"82004E40";
end if;
if pc = 21372 then
	inst <= x"07DC001C";
end if;
if pc = 21376 then
	inst <= x"8220538C";
end if;
if pc = 21380 then
	inst <= x"02200001";
end if;
if pc = 21384 then
	inst <= x"C1FDFFFC";
end if;
if pc = 21388 then
	inst <= x"C03C0010";
end if;
if pc = 21392 then
	inst <= x"02220001";
end if;
if pc = 21396 then
	inst <= x"22420220";
end if;
if pc = 21400 then
	inst <= x"C07C0004";
end if;
if pc = 21404 then
	inst <= x"D0464000";
end if;
if pc = 21408 then
	inst <= x"0280FFFF";
end if;
if pc = 21412 then
	inst <= x"824853F4";
end if;
if pc = 21416 then
	inst <= x"22440220";
end if;
if pc = 21420 then
	inst <= x"C09C0000";
end if;
if pc = 21424 then
	inst <= x"D0484000";
end if;
if pc = 21428 then
	inst <= x"02800000";
end if;
if pc = 21432 then
	inst <= x"C43C0014";
end if;
if pc = 21436 then
	inst <= x"C17DFFFC";
end if;
if pc = 21440 then
	inst <= x"00280000";
end if;
if pc = 21444 then
	inst <= x"03DC0020";
end if;
if pc = 21448 then
	inst <= x"037E000C";
end if;
if pc = 21452 then
	inst <= x"C57DFFFC";
end if;
if pc = 21456 then
	inst <= x"82004E40";
end if;
if pc = 21460 then
	inst <= x"07DC0020";
end if;
if pc = 21464 then
	inst <= x"822053E4";
end if;
if pc = 21468 then
	inst <= x"02200001";
end if;
if pc = 21472 then
	inst <= x"C1FDFFFC";
end if;
if pc = 21476 then
	inst <= x"C03C0014";
end if;
if pc = 21480 then
	inst <= x"02220001";
end if;
if pc = 21484 then
	inst <= x"C05C0004";
end if;
if pc = 21488 then
	inst <= x"82005284";
end if;
if pc = 21492 then
	inst <= x"02200000";
end if;
if pc = 21496 then
	inst <= x"C1FDFFFC";
end if;
if pc = 21500 then
	inst <= x"02200000";
end if;
if pc = 21504 then
	inst <= x"C1FDFFFC";
end if;
if pc = 21508 then
	inst <= x"02200000";
end if;
if pc = 21512 then
	inst <= x"C1FDFFFC";
end if;
if pc = 21516 then
	inst <= x"02200000";
end if;
if pc = 21520 then
	inst <= x"C1FDFFFC";
end if;
if pc = 21524 then
	inst <= x"22620220";
end if;
if pc = 21528 then
	inst <= x"D0646000";
end if;
if pc = 21532 then
	inst <= x"C0860000";
end if;
if pc = 21536 then
	inst <= x"02A0FFFF";
end if;
if pc = 21540 then
	inst <= x"828A57C0";
end if;
if pc = 21544 then
	inst <= x"02A00063";
end if;
if pc = 21548 then
	inst <= x"C47C0000";
end if;
if pc = 21552 then
	inst <= x"C45C0004";
end if;
if pc = 21556 then
	inst <= x"C43C0008";
end if;
if pc = 21560 then
	inst <= x"828A5678";
end if;
if pc = 21564 then
	inst <= x"02A00368";
end if;
if pc = 21568 then
	inst <= x"02C002B8";
end if;
if pc = 21572 then
	inst <= x"02E000C8";
end if;
if pc = 21576 then
	inst <= x"23080220";
end if;
if pc = 21580 then
	inst <= x"D0EF0000";
end if;
if pc = 21584 then
	inst <= x"C82C0000";
end if;
if pc = 21588 then
	inst <= x"C10E0014";
end if;
if pc = 21592 then
	inst <= x"C8500000";
end if;
if pc = 21596 then
	inst <= x"44224000";
end if;
if pc = 21600 then
	inst <= x"C84C0004";
end if;
if pc = 21604 then
	inst <= x"C10E0014";
end if;
if pc = 21608 then
	inst <= x"C8700004";
end if;
if pc = 21612 then
	inst <= x"44446000";
end if;
if pc = 21616 then
	inst <= x"C86C0008";
end if;
if pc = 21620 then
	inst <= x"C0CE0014";
end if;
if pc = 21624 then
	inst <= x"C88C0008";
end if;
if pc = 21628 then
	inst <= x"44668000";
end if;
if pc = 21632 then
	inst <= x"C0CA0004";
end if;
if pc = 21636 then
	inst <= x"22880220";
end if;
if pc = 21640 then
	inst <= x"D08C8000";
end if;
if pc = 21644 then
	inst <= x"C0CE0004";
end if;
if pc = 21648 then
	inst <= x"03000001";
end if;
if pc = 21652 then
	inst <= x"82D05504";
end if;
if pc = 21656 then
	inst <= x"02A00002";
end if;
if pc = 21660 then
	inst <= x"82CA54C4";
end if;
if pc = 21664 then
	inst <= x"C17DFFFC";
end if;
if pc = 21668 then
	inst <= x"00480000";
end if;
if pc = 21672 then
	inst <= x"002E0000";
end if;
if pc = 21676 then
	inst <= x"03DC0014";
end if;
if pc = 21680 then
	inst <= x"037E000C";
end if;
if pc = 21684 then
	inst <= x"C57DFFFC";
end if;
if pc = 21688 then
	inst <= x"82003A54";
end if;
if pc = 21692 then
	inst <= x"07DC0014";
end if;
if pc = 21696 then
	inst <= x"82005500";
end if;
if pc = 21700 then
	inst <= x"C8880000";
end if;
if pc = 21704 then
	inst <= x"8E8054D4";
end if;
if pc = 21708 then
	inst <= x"02200000";
end if;
if pc = 21712 then
	inst <= x"82005500";
end if;
if pc = 21716 then
	inst <= x"02A002AC";
end if;
if pc = 21720 then
	inst <= x"C8880004";
end if;
if pc = 21724 then
	inst <= x"48282000";
end if;
if pc = 21728 then
	inst <= x"C8880008";
end if;
if pc = 21732 then
	inst <= x"48484000";
end if;
if pc = 21736 then
	inst <= x"40224000";
end if;
if pc = 21740 then
	inst <= x"C848000C";
end if;
if pc = 21744 then
	inst <= x"48446000";
end if;
if pc = 21748 then
	inst <= x"40224000";
end if;
if pc = 21752 then
	inst <= x"CC2A0000";
end if;
if pc = 21756 then
	inst <= x"02200001";
end if;
if pc = 21760 then
	inst <= x"8200552C";
end if;
if pc = 21764 then
	inst <= x"C0AA0000";
end if;
if pc = 21768 then
	inst <= x"C17DFFFC";
end if;
if pc = 21772 then
	inst <= x"00680000";
end if;
if pc = 21776 then
	inst <= x"004A0000";
end if;
if pc = 21780 then
	inst <= x"002E0000";
end if;
if pc = 21784 then
	inst <= x"03DC0014";
end if;
if pc = 21788 then
	inst <= x"037E000C";
end if;
if pc = 21792 then
	inst <= x"C57DFFFC";
end if;
if pc = 21796 then
	inst <= x"8200389C";
end if;
if pc = 21800 then
	inst <= x"07DC0014";
end if;
if pc = 21804 then
	inst <= x"82205670";
end if;
if pc = 21808 then
	inst <= x"022002AC";
end if;
if pc = 21812 then
	inst <= x"C8220000";
end if;
if pc = 21816 then
	inst <= x"C8400070";
end if;
if pc = 21820 then
	inst <= x"8E245548";
end if;
if pc = 21824 then
	inst <= x"02200000";
end if;
if pc = 21828 then
	inst <= x"8200566C";
end if;
if pc = 21832 then
	inst <= x"C03C0000";
end if;
if pc = 21836 then
	inst <= x"C0420004";
end if;
if pc = 21840 then
	inst <= x"0260FFFF";
end if;
if pc = 21844 then
	inst <= x"82465658";
end if;
if pc = 21848 then
	inst <= x"026001E0";
end if;
if pc = 21852 then
	inst <= x"22440220";
end if;
if pc = 21856 then
	inst <= x"D0464000";
end if;
if pc = 21860 then
	inst <= x"02800000";
end if;
if pc = 21864 then
	inst <= x"C47C000C";
end if;
if pc = 21868 then
	inst <= x"C17DFFFC";
end if;
if pc = 21872 then
	inst <= x"00280000";
end if;
if pc = 21876 then
	inst <= x"03DC0018";
end if;
if pc = 21880 then
	inst <= x"037E000C";
end if;
if pc = 21884 then
	inst <= x"C57DFFFC";
end if;
if pc = 21888 then
	inst <= x"82004E40";
end if;
if pc = 21892 then
	inst <= x"07DC0018";
end if;
if pc = 21896 then
	inst <= x"82205594";
end if;
if pc = 21900 then
	inst <= x"02200001";
end if;
if pc = 21904 then
	inst <= x"82005654";
end if;
if pc = 21908 then
	inst <= x"C03C0000";
end if;
if pc = 21912 then
	inst <= x"C0420008";
end if;
if pc = 21916 then
	inst <= x"0260FFFF";
end if;
if pc = 21920 then
	inst <= x"82465650";
end if;
if pc = 21924 then
	inst <= x"22440220";
end if;
if pc = 21928 then
	inst <= x"C07C000C";
end if;
if pc = 21932 then
	inst <= x"D0464000";
end if;
if pc = 21936 then
	inst <= x"02800000";
end if;
if pc = 21940 then
	inst <= x"C17DFFFC";
end if;
if pc = 21944 then
	inst <= x"00280000";
end if;
if pc = 21948 then
	inst <= x"03DC0018";
end if;
if pc = 21952 then
	inst <= x"037E000C";
end if;
if pc = 21956 then
	inst <= x"C57DFFFC";
end if;
if pc = 21960 then
	inst <= x"82004E40";
end if;
if pc = 21964 then
	inst <= x"07DC0018";
end if;
if pc = 21968 then
	inst <= x"822055DC";
end if;
if pc = 21972 then
	inst <= x"02200001";
end if;
if pc = 21976 then
	inst <= x"8200564C";
end if;
if pc = 21980 then
	inst <= x"C03C0000";
end if;
if pc = 21984 then
	inst <= x"C042000C";
end if;
if pc = 21988 then
	inst <= x"0260FFFF";
end if;
if pc = 21992 then
	inst <= x"82465648";
end if;
if pc = 21996 then
	inst <= x"22440220";
end if;
if pc = 22000 then
	inst <= x"C07C000C";
end if;
if pc = 22004 then
	inst <= x"D0464000";
end if;
if pc = 22008 then
	inst <= x"02600000";
end if;
if pc = 22012 then
	inst <= x"C17DFFFC";
end if;
if pc = 22016 then
	inst <= x"00260000";
end if;
if pc = 22020 then
	inst <= x"03DC0018";
end if;
if pc = 22024 then
	inst <= x"037E000C";
end if;
if pc = 22028 then
	inst <= x"C57DFFFC";
end if;
if pc = 22032 then
	inst <= x"82004E40";
end if;
if pc = 22036 then
	inst <= x"07DC0018";
end if;
if pc = 22040 then
	inst <= x"82205624";
end if;
if pc = 22044 then
	inst <= x"02200001";
end if;
if pc = 22048 then
	inst <= x"82005644";
end if;
if pc = 22052 then
	inst <= x"02200004";
end if;
if pc = 22056 then
	inst <= x"C05C0000";
end if;
if pc = 22060 then
	inst <= x"C17DFFFC";
end if;
if pc = 22064 then
	inst <= x"03DC0018";
end if;
if pc = 22068 then
	inst <= x"037E000C";
end if;
if pc = 22072 then
	inst <= x"C57DFFFC";
end if;
if pc = 22076 then
	inst <= x"82005284";
end if;
if pc = 22080 then
	inst <= x"07DC0018";
end if;
if pc = 22084 then
	inst <= x"8200564C";
end if;
if pc = 22088 then
	inst <= x"02200000";
end if;
if pc = 22092 then
	inst <= x"82005654";
end if;
if pc = 22096 then
	inst <= x"02200000";
end if;
if pc = 22100 then
	inst <= x"8200565C";
end if;
if pc = 22104 then
	inst <= x"02200000";
end if;
if pc = 22108 then
	inst <= x"82205668";
end if;
if pc = 22112 then
	inst <= x"02200001";
end if;
if pc = 22116 then
	inst <= x"8200566C";
end if;
if pc = 22120 then
	inst <= x"02200000";
end if;
if pc = 22124 then
	inst <= x"82005674";
end if;
if pc = 22128 then
	inst <= x"02200000";
end if;
if pc = 22132 then
	inst <= x"8200567C";
end if;
if pc = 22136 then
	inst <= x"02200001";
end if;
if pc = 22140 then
	inst <= x"822057B0";
end if;
if pc = 22144 then
	inst <= x"C03C0000";
end if;
if pc = 22148 then
	inst <= x"C0420004";
end if;
if pc = 22152 then
	inst <= x"0260FFFF";
end if;
if pc = 22156 then
	inst <= x"82465790";
end if;
if pc = 22160 then
	inst <= x"026001E0";
end if;
if pc = 22164 then
	inst <= x"22440220";
end if;
if pc = 22168 then
	inst <= x"D0464000";
end if;
if pc = 22172 then
	inst <= x"02800000";
end if;
if pc = 22176 then
	inst <= x"C47C0010";
end if;
if pc = 22180 then
	inst <= x"C17DFFFC";
end if;
if pc = 22184 then
	inst <= x"00280000";
end if;
if pc = 22188 then
	inst <= x"03DC001C";
end if;
if pc = 22192 then
	inst <= x"037E000C";
end if;
if pc = 22196 then
	inst <= x"C57DFFFC";
end if;
if pc = 22200 then
	inst <= x"82004E40";
end if;
if pc = 22204 then
	inst <= x"07DC001C";
end if;
if pc = 22208 then
	inst <= x"822056CC";
end if;
if pc = 22212 then
	inst <= x"02200001";
end if;
if pc = 22216 then
	inst <= x"8200578C";
end if;
if pc = 22220 then
	inst <= x"C03C0000";
end if;
if pc = 22224 then
	inst <= x"C0420008";
end if;
if pc = 22228 then
	inst <= x"0260FFFF";
end if;
if pc = 22232 then
	inst <= x"82465788";
end if;
if pc = 22236 then
	inst <= x"22440220";
end if;
if pc = 22240 then
	inst <= x"C07C0010";
end if;
if pc = 22244 then
	inst <= x"D0464000";
end if;
if pc = 22248 then
	inst <= x"02800000";
end if;
if pc = 22252 then
	inst <= x"C17DFFFC";
end if;
if pc = 22256 then
	inst <= x"00280000";
end if;
if pc = 22260 then
	inst <= x"03DC001C";
end if;
if pc = 22264 then
	inst <= x"037E000C";
end if;
if pc = 22268 then
	inst <= x"C57DFFFC";
end if;
if pc = 22272 then
	inst <= x"82004E40";
end if;
if pc = 22276 then
	inst <= x"07DC001C";
end if;
if pc = 22280 then
	inst <= x"82205714";
end if;
if pc = 22284 then
	inst <= x"02200001";
end if;
if pc = 22288 then
	inst <= x"82005784";
end if;
if pc = 22292 then
	inst <= x"C03C0000";
end if;
if pc = 22296 then
	inst <= x"C042000C";
end if;
if pc = 22300 then
	inst <= x"0260FFFF";
end if;
if pc = 22304 then
	inst <= x"82465780";
end if;
if pc = 22308 then
	inst <= x"22440220";
end if;
if pc = 22312 then
	inst <= x"C07C0010";
end if;
if pc = 22316 then
	inst <= x"D0464000";
end if;
if pc = 22320 then
	inst <= x"02600000";
end if;
if pc = 22324 then
	inst <= x"C17DFFFC";
end if;
if pc = 22328 then
	inst <= x"00260000";
end if;
if pc = 22332 then
	inst <= x"03DC001C";
end if;
if pc = 22336 then
	inst <= x"037E000C";
end if;
if pc = 22340 then
	inst <= x"C57DFFFC";
end if;
if pc = 22344 then
	inst <= x"82004E40";
end if;
if pc = 22348 then
	inst <= x"07DC001C";
end if;
if pc = 22352 then
	inst <= x"8220575C";
end if;
if pc = 22356 then
	inst <= x"02200001";
end if;
if pc = 22360 then
	inst <= x"8200577C";
end if;
if pc = 22364 then
	inst <= x"02200004";
end if;
if pc = 22368 then
	inst <= x"C05C0000";
end if;
if pc = 22372 then
	inst <= x"C17DFFFC";
end if;
if pc = 22376 then
	inst <= x"03DC001C";
end if;
if pc = 22380 then
	inst <= x"037E000C";
end if;
if pc = 22384 then
	inst <= x"C57DFFFC";
end if;
if pc = 22388 then
	inst <= x"82005284";
end if;
if pc = 22392 then
	inst <= x"07DC001C";
end if;
if pc = 22396 then
	inst <= x"82005784";
end if;
if pc = 22400 then
	inst <= x"02200000";
end if;
if pc = 22404 then
	inst <= x"8200578C";
end if;
if pc = 22408 then
	inst <= x"02200000";
end if;
if pc = 22412 then
	inst <= x"82005794";
end if;
if pc = 22416 then
	inst <= x"02200000";
end if;
if pc = 22420 then
	inst <= x"822057A0";
end if;
if pc = 22424 then
	inst <= x"02200001";
end if;
if pc = 22428 then
	inst <= x"C1FDFFFC";
end if;
if pc = 22432 then
	inst <= x"C03C0008";
end if;
if pc = 22436 then
	inst <= x"02220001";
end if;
if pc = 22440 then
	inst <= x"C05C0004";
end if;
if pc = 22444 then
	inst <= x"82005414";
end if;
if pc = 22448 then
	inst <= x"C03C0008";
end if;
if pc = 22452 then
	inst <= x"02220001";
end if;
if pc = 22456 then
	inst <= x"C05C0004";
end if;
if pc = 22460 then
	inst <= x"82005414";
end if;
if pc = 22464 then
	inst <= x"02200000";
end if;
if pc = 22468 then
	inst <= x"C1FDFFFC";
end if;
if pc = 22472 then
	inst <= x"22820220";
end if;
if pc = 22476 then
	inst <= x"D0848000";
end if;
if pc = 22480 then
	inst <= x"02A0FFFF";
end if;
if pc = 22484 then
	inst <= x"828A5CD8";
end if;
if pc = 22488 then
	inst <= x"02A0030C";
end if;
if pc = 22492 then
	inst <= x"02C000C8";
end if;
if pc = 22496 then
	inst <= x"22E80220";
end if;
if pc = 22500 then
	inst <= x"D0ECE000";
end if;
if pc = 22504 then
	inst <= x"C82A0000";
end if;
if pc = 22508 then
	inst <= x"C10E0014";
end if;
if pc = 22512 then
	inst <= x"C8500000";
end if;
if pc = 22516 then
	inst <= x"44224000";
end if;
if pc = 22520 then
	inst <= x"C84A0004";
end if;
if pc = 22524 then
	inst <= x"C10E0014";
end if;
if pc = 22528 then
	inst <= x"C8700004";
end if;
if pc = 22532 then
	inst <= x"44446000";
end if;
if pc = 22536 then
	inst <= x"C86A0008";
end if;
if pc = 22540 then
	inst <= x"C10E0014";
end if;
if pc = 22544 then
	inst <= x"C8900008";
end if;
if pc = 22548 then
	inst <= x"44668000";
end if;
if pc = 22552 then
	inst <= x"C10E0004";
end if;
if pc = 22556 then
	inst <= x"03200001";
end if;
if pc = 22560 then
	inst <= x"C4BC0000";
end if;
if pc = 22564 then
	inst <= x"C47C0004";
end if;
if pc = 22568 then
	inst <= x"C45C0008";
end if;
if pc = 22572 then
	inst <= x"C43C000C";
end if;
if pc = 22576 then
	inst <= x"C4DC0010";
end if;
if pc = 22580 then
	inst <= x"C49C0014";
end if;
if pc = 22584 then
	inst <= x"8312588C";
end if;
if pc = 22588 then
	inst <= x"03200002";
end if;
if pc = 22592 then
	inst <= x"83125868";
end if;
if pc = 22596 then
	inst <= x"C17DFFFC";
end if;
if pc = 22600 then
	inst <= x"00460000";
end if;
if pc = 22604 then
	inst <= x"002E0000";
end if;
if pc = 22608 then
	inst <= x"03DC0020";
end if;
if pc = 22612 then
	inst <= x"037E000C";
end if;
if pc = 22616 then
	inst <= x"C57DFFFC";
end if;
if pc = 22620 then
	inst <= x"820034A0";
end if;
if pc = 22624 then
	inst <= x"07DC0020";
end if;
if pc = 22628 then
	inst <= x"82005888";
end if;
if pc = 22632 then
	inst <= x"C17DFFFC";
end if;
if pc = 22636 then
	inst <= x"00460000";
end if;
if pc = 22640 then
	inst <= x"002E0000";
end if;
if pc = 22644 then
	inst <= x"03DC0020";
end if;
if pc = 22648 then
	inst <= x"037E000C";
end if;
if pc = 22652 then
	inst <= x"C57DFFFC";
end if;
if pc = 22656 then
	inst <= x"820032A4";
end if;
if pc = 22660 then
	inst <= x"07DC0020";
end if;
if pc = 22664 then
	inst <= x"8200596C";
end if;
if pc = 22668 then
	inst <= x"03000000";
end if;
if pc = 22672 then
	inst <= x"03200001";
end if;
if pc = 22676 then
	inst <= x"03400002";
end if;
if pc = 22680 then
	inst <= x"CC3C0018";
end if;
if pc = 22684 then
	inst <= x"CC7C0020";
end if;
if pc = 22688 then
	inst <= x"CC5C0028";
end if;
if pc = 22692 then
	inst <= x"C4FC0030";
end if;
if pc = 22696 then
	inst <= x"C17DFFFC";
end if;
if pc = 22700 then
	inst <= x"00B40000";
end if;
if pc = 22704 then
	inst <= x"00920000";
end if;
if pc = 22708 then
	inst <= x"00460000";
end if;
if pc = 22712 then
	inst <= x"002E0000";
end if;
if pc = 22716 then
	inst <= x"00700000";
end if;
if pc = 22720 then
	inst <= x"03DC003C";
end if;
if pc = 22724 then
	inst <= x"037E000C";
end if;
if pc = 22728 then
	inst <= x"C57DFFFC";
end if;
if pc = 22732 then
	inst <= x"8200317C";
end if;
if pc = 22736 then
	inst <= x"07DC003C";
end if;
if pc = 22740 then
	inst <= x"822058E0";
end if;
if pc = 22744 then
	inst <= x"02200001";
end if;
if pc = 22748 then
	inst <= x"8200596C";
end if;
if pc = 22752 then
	inst <= x"02600001";
end if;
if pc = 22756 then
	inst <= x"02800002";
end if;
if pc = 22760 then
	inst <= x"02A00000";
end if;
if pc = 22764 then
	inst <= x"C83C0028";
end if;
if pc = 22768 then
	inst <= x"C85C0020";
end if;
if pc = 22772 then
	inst <= x"C87C0018";
end if;
if pc = 22776 then
	inst <= x"C03C0030";
end if;
if pc = 22780 then
	inst <= x"C05C0004";
end if;
if pc = 22784 then
	inst <= x"C17DFFFC";
end if;
if pc = 22788 then
	inst <= x"03DC003C";
end if;
if pc = 22792 then
	inst <= x"037E000C";
end if;
if pc = 22796 then
	inst <= x"C57DFFFC";
end if;
if pc = 22800 then
	inst <= x"8200317C";
end if;
if pc = 22804 then
	inst <= x"07DC003C";
end if;
if pc = 22808 then
	inst <= x"82205924";
end if;
if pc = 22812 then
	inst <= x"02200002";
end if;
if pc = 22816 then
	inst <= x"8200596C";
end if;
if pc = 22820 then
	inst <= x"02600002";
end if;
if pc = 22824 then
	inst <= x"02800000";
end if;
if pc = 22828 then
	inst <= x"02A00001";
end if;
if pc = 22832 then
	inst <= x"C83C0020";
end if;
if pc = 22836 then
	inst <= x"C85C0018";
end if;
if pc = 22840 then
	inst <= x"C87C0028";
end if;
if pc = 22844 then
	inst <= x"C03C0030";
end if;
if pc = 22848 then
	inst <= x"C05C0004";
end if;
if pc = 22852 then
	inst <= x"C17DFFFC";
end if;
if pc = 22856 then
	inst <= x"03DC003C";
end if;
if pc = 22860 then
	inst <= x"037E000C";
end if;
if pc = 22864 then
	inst <= x"C57DFFFC";
end if;
if pc = 22868 then
	inst <= x"8200317C";
end if;
if pc = 22872 then
	inst <= x"07DC003C";
end if;
if pc = 22876 then
	inst <= x"82205968";
end if;
if pc = 22880 then
	inst <= x"02200003";
end if;
if pc = 22884 then
	inst <= x"8200596C";
end if;
if pc = 22888 then
	inst <= x"02200000";
end if;
if pc = 22892 then
	inst <= x"82205CA8";
end if;
if pc = 22896 then
	inst <= x"024002AC";
end if;
if pc = 22900 then
	inst <= x"C8240000";
end if;
if pc = 22904 then
	inst <= x"8E025980";
end if;
if pc = 22908 then
	inst <= x"82005C94";
end if;
if pc = 22912 then
	inst <= x"024002B4";
end if;
if pc = 22916 then
	inst <= x"C8440000";
end if;
if pc = 22920 then
	inst <= x"8E245990";
end if;
if pc = 22924 then
	inst <= x"82005C94";
end if;
if pc = 22928 then
	inst <= x"C8400074";
end if;
if pc = 22932 then
	inst <= x"40224000";
end if;
if pc = 22936 then
	inst <= x"C07C0004";
end if;
if pc = 22940 then
	inst <= x"C8460000";
end if;
if pc = 22944 then
	inst <= x"48442000";
end if;
if pc = 22948 then
	inst <= x"C09C0000";
end if;
if pc = 22952 then
	inst <= x"C8680000";
end if;
if pc = 22956 then
	inst <= x"40446000";
end if;
if pc = 22960 then
	inst <= x"C8660004";
end if;
if pc = 22964 then
	inst <= x"48662000";
end if;
if pc = 22968 then
	inst <= x"C8880004";
end if;
if pc = 22972 then
	inst <= x"40668000";
end if;
if pc = 22976 then
	inst <= x"C8860008";
end if;
if pc = 22980 then
	inst <= x"48882000";
end if;
if pc = 22984 then
	inst <= x"C8A80008";
end if;
if pc = 22988 then
	inst <= x"4088A000";
end if;
if pc = 22992 then
	inst <= x"C09C0008";
end if;
if pc = 22996 then
	inst <= x"C0A80000";
end if;
if pc = 23000 then
	inst <= x"02C0FFFF";
end if;
if pc = 23004 then
	inst <= x"C43C0034";
end if;
if pc = 23008 then
	inst <= x"CC9C0038";
end if;
if pc = 23012 then
	inst <= x"CC7C0040";
end if;
if pc = 23016 then
	inst <= x"CC5C0048";
end if;
if pc = 23020 then
	inst <= x"C45C0050";
end if;
if pc = 23024 then
	inst <= x"CC3C0058";
end if;
if pc = 23028 then
	inst <= x"82AC5C48";
end if;
if pc = 23032 then
	inst <= x"22AA0220";
end if;
if pc = 23036 then
	inst <= x"C0DC0010";
end if;
if pc = 23040 then
	inst <= x"D0ACA000";
end if;
if pc = 23044 then
	inst <= x"C17DFFFC";
end if;
if pc = 23048 then
	inst <= x"002A0000";
end if;
if pc = 23052 then
	inst <= x"40204000";
end if;
if pc = 23056 then
	inst <= x"40406000";
end if;
if pc = 23060 then
	inst <= x"40608000";
end if;
if pc = 23064 then
	inst <= x"03DC0068";
end if;
if pc = 23068 then
	inst <= x"037E000C";
end if;
if pc = 23072 then
	inst <= x"C57DFFFC";
end if;
if pc = 23076 then
	inst <= x"82004860";
end if;
if pc = 23080 then
	inst <= x"07DC0068";
end if;
if pc = 23084 then
	inst <= x"82205A38";
end if;
if pc = 23088 then
	inst <= x"02200000";
end if;
if pc = 23092 then
	inst <= x"82005C44";
end if;
if pc = 23096 then
	inst <= x"C05C0008";
end if;
if pc = 23100 then
	inst <= x"C0240004";
end if;
if pc = 23104 then
	inst <= x"0260FFFF";
end if;
if pc = 23108 then
	inst <= x"82265C40";
end if;
if pc = 23112 then
	inst <= x"22220220";
end if;
if pc = 23116 then
	inst <= x"C07C0010";
end if;
if pc = 23120 then
	inst <= x"D0262000";
end if;
if pc = 23124 then
	inst <= x"C0820014";
end if;
if pc = 23128 then
	inst <= x"C8280000";
end if;
if pc = 23132 then
	inst <= x"C85C0048";
end if;
if pc = 23136 then
	inst <= x"44242000";
end if;
if pc = 23140 then
	inst <= x"C0820014";
end if;
if pc = 23144 then
	inst <= x"C8680004";
end if;
if pc = 23148 then
	inst <= x"C89C0040";
end if;
if pc = 23152 then
	inst <= x"44686000";
end if;
if pc = 23156 then
	inst <= x"C0820014";
end if;
if pc = 23160 then
	inst <= x"C8A80008";
end if;
if pc = 23164 then
	inst <= x"C8DC0038";
end if;
if pc = 23168 then
	inst <= x"44ACA000";
end if;
if pc = 23172 then
	inst <= x"C0820004";
end if;
if pc = 23176 then
	inst <= x"02A00001";
end if;
if pc = 23180 then
	inst <= x"828A5B24";
end if;
if pc = 23184 then
	inst <= x"02A00002";
end if;
if pc = 23188 then
	inst <= x"828A5ABC";
end if;
if pc = 23192 then
	inst <= x"C17DFFFC";
end if;
if pc = 23196 then
	inst <= x"40406000";
end if;
if pc = 23200 then
	inst <= x"4060A000";
end if;
if pc = 23204 then
	inst <= x"03DC0068";
end if;
if pc = 23208 then
	inst <= x"037E000C";
end if;
if pc = 23212 then
	inst <= x"C57DFFFC";
end if;
if pc = 23216 then
	inst <= x"82004780";
end if;
if pc = 23220 then
	inst <= x"07DC0068";
end if;
if pc = 23224 then
	inst <= x"82005B20";
end if;
if pc = 23228 then
	inst <= x"C0820010";
end if;
if pc = 23232 then
	inst <= x"C8E80000";
end if;
if pc = 23236 then
	inst <= x"482E2000";
end if;
if pc = 23240 then
	inst <= x"C8E80004";
end if;
if pc = 23244 then
	inst <= x"486E6000";
end if;
if pc = 23248 then
	inst <= x"40226000";
end if;
if pc = 23252 then
	inst <= x"C8680008";
end if;
if pc = 23256 then
	inst <= x"4866A000";
end if;
if pc = 23260 then
	inst <= x"40226000";
end if;
if pc = 23264 then
	inst <= x"C0220018";
end if;
if pc = 23268 then
	inst <= x"8E205AF0";
end if;
if pc = 23272 then
	inst <= x"02800000";
end if;
if pc = 23276 then
	inst <= x"82005AF4";
end if;
if pc = 23280 then
	inst <= x"02800001";
end if;
if pc = 23284 then
	inst <= x"82205B0C";
end if;
if pc = 23288 then
	inst <= x"8E205B04";
end if;
if pc = 23292 then
	inst <= x"02200001";
end if;
if pc = 23296 then
	inst <= x"82005B08";
end if;
if pc = 23300 then
	inst <= x"02200000";
end if;
if pc = 23304 then
	inst <= x"82005B10";
end if;
if pc = 23308 then
	inst <= x"00280000";
end if;
if pc = 23312 then
	inst <= x"82205B1C";
end if;
if pc = 23316 then
	inst <= x"02200000";
end if;
if pc = 23320 then
	inst <= x"82005B20";
end if;
if pc = 23324 then
	inst <= x"02200001";
end if;
if pc = 23328 then
	inst <= x"82005BB0";
end if;
if pc = 23332 then
	inst <= x"8E205B2C";
end if;
if pc = 23336 then
	inst <= x"82005B30";
end if;
if pc = 23340 then
	inst <= x"44202000";
end if;
if pc = 23344 then
	inst <= x"C0820010";
end if;
if pc = 23348 then
	inst <= x"C8E80000";
end if;
if pc = 23352 then
	inst <= x"8E2E5B44";
end if;
if pc = 23356 then
	inst <= x"02800000";
end if;
if pc = 23360 then
	inst <= x"82005B90";
end if;
if pc = 23364 then
	inst <= x"8E605B50";
end if;
if pc = 23368 then
	inst <= x"40206000";
end if;
if pc = 23372 then
	inst <= x"82005B54";
end if;
if pc = 23376 then
	inst <= x"44206000";
end if;
if pc = 23380 then
	inst <= x"C0820010";
end if;
if pc = 23384 then
	inst <= x"C8680004";
end if;
if pc = 23388 then
	inst <= x"8E265B68";
end if;
if pc = 23392 then
	inst <= x"02800000";
end if;
if pc = 23396 then
	inst <= x"82005B90";
end if;
if pc = 23400 then
	inst <= x"8EA05B74";
end if;
if pc = 23404 then
	inst <= x"4020A000";
end if;
if pc = 23408 then
	inst <= x"82005B78";
end if;
if pc = 23412 then
	inst <= x"4420A000";
end if;
if pc = 23416 then
	inst <= x"C0820010";
end if;
if pc = 23420 then
	inst <= x"C8680008";
end if;
if pc = 23424 then
	inst <= x"8E265B8C";
end if;
if pc = 23428 then
	inst <= x"02800000";
end if;
if pc = 23432 then
	inst <= x"82005B90";
end if;
if pc = 23436 then
	inst <= x"02800001";
end if;
if pc = 23440 then
	inst <= x"82805B9C";
end if;
if pc = 23444 then
	inst <= x"C0220018";
end if;
if pc = 23448 then
	inst <= x"82005BB0";
end if;
if pc = 23452 then
	inst <= x"C0220018";
end if;
if pc = 23456 then
	inst <= x"82205BAC";
end if;
if pc = 23460 then
	inst <= x"02200000";
end if;
if pc = 23464 then
	inst <= x"82005BB0";
end if;
if pc = 23468 then
	inst <= x"02200001";
end if;
if pc = 23472 then
	inst <= x"82205BBC";
end if;
if pc = 23476 then
	inst <= x"02200000";
end if;
if pc = 23480 then
	inst <= x"82005C3C";
end if;
if pc = 23484 then
	inst <= x"C05C0008";
end if;
if pc = 23488 then
	inst <= x"C0240008";
end if;
if pc = 23492 then
	inst <= x"0260FFFF";
end if;
if pc = 23496 then
	inst <= x"82265C38";
end if;
if pc = 23500 then
	inst <= x"22220220";
end if;
if pc = 23504 then
	inst <= x"C07C0010";
end if;
if pc = 23508 then
	inst <= x"D0262000";
end if;
if pc = 23512 then
	inst <= x"C83C0048";
end if;
if pc = 23516 then
	inst <= x"C85C0040";
end if;
if pc = 23520 then
	inst <= x"C87C0038";
end if;
if pc = 23524 then
	inst <= x"C17DFFFC";
end if;
if pc = 23528 then
	inst <= x"03DC0068";
end if;
if pc = 23532 then
	inst <= x"037E000C";
end if;
if pc = 23536 then
	inst <= x"C57DFFFC";
end if;
if pc = 23540 then
	inst <= x"82004860";
end if;
if pc = 23544 then
	inst <= x"07DC0068";
end if;
if pc = 23548 then
	inst <= x"82205C08";
end if;
if pc = 23552 then
	inst <= x"02200000";
end if;
if pc = 23556 then
	inst <= x"82005C34";
end if;
if pc = 23560 then
	inst <= x"02200003";
end if;
if pc = 23564 then
	inst <= x"C83C0048";
end if;
if pc = 23568 then
	inst <= x"C85C0040";
end if;
if pc = 23572 then
	inst <= x"C87C0038";
end if;
if pc = 23576 then
	inst <= x"C05C0008";
end if;
if pc = 23580 then
	inst <= x"C17DFFFC";
end if;
if pc = 23584 then
	inst <= x"03DC0068";
end if;
if pc = 23588 then
	inst <= x"037E000C";
end if;
if pc = 23592 then
	inst <= x"C57DFFFC";
end if;
if pc = 23596 then
	inst <= x"82004A0C";
end if;
if pc = 23600 then
	inst <= x"07DC0068";
end if;
if pc = 23604 then
	inst <= x"82005C3C";
end if;
if pc = 23608 then
	inst <= x"02200001";
end if;
if pc = 23612 then
	inst <= x"82005C44";
end if;
if pc = 23616 then
	inst <= x"02200001";
end if;
if pc = 23620 then
	inst <= x"82005C4C";
end if;
if pc = 23624 then
	inst <= x"02200001";
end if;
if pc = 23628 then
	inst <= x"82205C94";
end if;
if pc = 23632 then
	inst <= x"C03C0050";
end if;
if pc = 23636 then
	inst <= x"C83C0058";
end if;
if pc = 23640 then
	inst <= x"CC220000";
end if;
if pc = 23644 then
	inst <= x"022002B8";
end if;
if pc = 23648 then
	inst <= x"C83C0048";
end if;
if pc = 23652 then
	inst <= x"CC220000";
end if;
if pc = 23656 then
	inst <= x"C83C0040";
end if;
if pc = 23660 then
	inst <= x"CC220004";
end if;
if pc = 23664 then
	inst <= x"C83C0038";
end if;
if pc = 23668 then
	inst <= x"CC220008";
end if;
if pc = 23672 then
	inst <= x"022002C4";
end if;
if pc = 23676 then
	inst <= x"C05C0014";
end if;
if pc = 23680 then
	inst <= x"C4420000";
end if;
if pc = 23684 then
	inst <= x"022002B0";
end if;
if pc = 23688 then
	inst <= x"C05C0034";
end if;
if pc = 23692 then
	inst <= x"C4420000";
end if;
if pc = 23696 then
	inst <= x"82005C94";
end if;
if pc = 23700 then
	inst <= x"C03C000C";
end if;
if pc = 23704 then
	inst <= x"02220001";
end if;
if pc = 23708 then
	inst <= x"C05C0008";
end if;
if pc = 23712 then
	inst <= x"C07C0004";
end if;
if pc = 23716 then
	inst <= x"820057C8";
end if;
if pc = 23720 then
	inst <= x"C03C0014";
end if;
if pc = 23724 then
	inst <= x"22220220";
end if;
if pc = 23728 then
	inst <= x"C05C0010";
end if;
if pc = 23732 then
	inst <= x"D0242000";
end if;
if pc = 23736 then
	inst <= x"C0220018";
end if;
if pc = 23740 then
	inst <= x"82205CD4";
end if;
if pc = 23744 then
	inst <= x"C03C000C";
end if;
if pc = 23748 then
	inst <= x"02220001";
end if;
if pc = 23752 then
	inst <= x"C05C0008";
end if;
if pc = 23756 then
	inst <= x"C07C0004";
end if;
if pc = 23760 then
	inst <= x"820057C8";
end if;
if pc = 23764 then
	inst <= x"C1FDFFFC";
end if;
if pc = 23768 then
	inst <= x"C1FDFFFC";
end if;
if pc = 23772 then
	inst <= x"22820220";
end if;
if pc = 23776 then
	inst <= x"D0848000";
end if;
if pc = 23780 then
	inst <= x"02A0FFFF";
end if;
if pc = 23784 then
	inst <= x"828A5E48";
end if;
if pc = 23788 then
	inst <= x"02A001E0";
end if;
if pc = 23792 then
	inst <= x"22880220";
end if;
if pc = 23796 then
	inst <= x"D08A8000";
end if;
if pc = 23800 then
	inst <= x"02C00000";
end if;
if pc = 23804 then
	inst <= x"C47C0000";
end if;
if pc = 23808 then
	inst <= x"C4BC0004";
end if;
if pc = 23812 then
	inst <= x"C45C0008";
end if;
if pc = 23816 then
	inst <= x"C43C000C";
end if;
if pc = 23820 then
	inst <= x"C17DFFFC";
end if;
if pc = 23824 then
	inst <= x"00480000";
end if;
if pc = 23828 then
	inst <= x"002C0000";
end if;
if pc = 23832 then
	inst <= x"03DC0018";
end if;
if pc = 23836 then
	inst <= x"037E000C";
end if;
if pc = 23840 then
	inst <= x"C57DFFFC";
end if;
if pc = 23844 then
	inst <= x"820057C8";
end if;
if pc = 23848 then
	inst <= x"07DC0018";
end if;
if pc = 23852 then
	inst <= x"C03C000C";
end if;
if pc = 23856 then
	inst <= x"02220001";
end if;
if pc = 23860 then
	inst <= x"22420220";
end if;
if pc = 23864 then
	inst <= x"C07C0008";
end if;
if pc = 23868 then
	inst <= x"D0464000";
end if;
if pc = 23872 then
	inst <= x"0280FFFF";
end if;
if pc = 23876 then
	inst <= x"82485E44";
end if;
if pc = 23880 then
	inst <= x"22440220";
end if;
if pc = 23884 then
	inst <= x"C09C0004";
end if;
if pc = 23888 then
	inst <= x"D0484000";
end if;
if pc = 23892 then
	inst <= x"02A00000";
end if;
if pc = 23896 then
	inst <= x"C0DC0000";
end if;
if pc = 23900 then
	inst <= x"C43C0010";
end if;
if pc = 23904 then
	inst <= x"C17DFFFC";
end if;
if pc = 23908 then
	inst <= x"006C0000";
end if;
if pc = 23912 then
	inst <= x"002A0000";
end if;
if pc = 23916 then
	inst <= x"03DC001C";
end if;
if pc = 23920 then
	inst <= x"037E000C";
end if;
if pc = 23924 then
	inst <= x"C57DFFFC";
end if;
if pc = 23928 then
	inst <= x"820057C8";
end if;
if pc = 23932 then
	inst <= x"07DC001C";
end if;
if pc = 23936 then
	inst <= x"C03C0010";
end if;
if pc = 23940 then
	inst <= x"02220001";
end if;
if pc = 23944 then
	inst <= x"22420220";
end if;
if pc = 23948 then
	inst <= x"C07C0008";
end if;
if pc = 23952 then
	inst <= x"D0464000";
end if;
if pc = 23956 then
	inst <= x"0280FFFF";
end if;
if pc = 23960 then
	inst <= x"82485E40";
end if;
if pc = 23964 then
	inst <= x"22440220";
end if;
if pc = 23968 then
	inst <= x"C09C0004";
end if;
if pc = 23972 then
	inst <= x"D0484000";
end if;
if pc = 23976 then
	inst <= x"02A00000";
end if;
if pc = 23980 then
	inst <= x"C0DC0000";
end if;
if pc = 23984 then
	inst <= x"C43C0014";
end if;
if pc = 23988 then
	inst <= x"C17DFFFC";
end if;
if pc = 23992 then
	inst <= x"006C0000";
end if;
if pc = 23996 then
	inst <= x"002A0000";
end if;
if pc = 24000 then
	inst <= x"03DC0020";
end if;
if pc = 24004 then
	inst <= x"037E000C";
end if;
if pc = 24008 then
	inst <= x"C57DFFFC";
end if;
if pc = 24012 then
	inst <= x"820057C8";
end if;
if pc = 24016 then
	inst <= x"07DC0020";
end if;
if pc = 24020 then
	inst <= x"C03C0014";
end if;
if pc = 24024 then
	inst <= x"02220001";
end if;
if pc = 24028 then
	inst <= x"22420220";
end if;
if pc = 24032 then
	inst <= x"C07C0008";
end if;
if pc = 24036 then
	inst <= x"D0464000";
end if;
if pc = 24040 then
	inst <= x"0280FFFF";
end if;
if pc = 24044 then
	inst <= x"82485E3C";
end if;
if pc = 24048 then
	inst <= x"22440220";
end if;
if pc = 24052 then
	inst <= x"C09C0004";
end if;
if pc = 24056 then
	inst <= x"D0484000";
end if;
if pc = 24060 then
	inst <= x"02800000";
end if;
if pc = 24064 then
	inst <= x"C0BC0000";
end if;
if pc = 24068 then
	inst <= x"C43C0018";
end if;
if pc = 24072 then
	inst <= x"C17DFFFC";
end if;
if pc = 24076 then
	inst <= x"006A0000";
end if;
if pc = 24080 then
	inst <= x"00280000";
end if;
if pc = 24084 then
	inst <= x"03DC0024";
end if;
if pc = 24088 then
	inst <= x"037E000C";
end if;
if pc = 24092 then
	inst <= x"C57DFFFC";
end if;
if pc = 24096 then
	inst <= x"820057C8";
end if;
if pc = 24100 then
	inst <= x"07DC0024";
end if;
if pc = 24104 then
	inst <= x"C03C0018";
end if;
if pc = 24108 then
	inst <= x"02220001";
end if;
if pc = 24112 then
	inst <= x"C05C0008";
end if;
if pc = 24116 then
	inst <= x"C07C0000";
end if;
if pc = 24120 then
	inst <= x"82005CDC";
end if;
if pc = 24124 then
	inst <= x"C1FDFFFC";
end if;
if pc = 24128 then
	inst <= x"C1FDFFFC";
end if;
if pc = 24132 then
	inst <= x"C1FDFFFC";
end if;
if pc = 24136 then
	inst <= x"C1FDFFFC";
end if;
if pc = 24140 then
	inst <= x"22820220";
end if;
if pc = 24144 then
	inst <= x"D0848000";
end if;
if pc = 24148 then
	inst <= x"C0A80000";
end if;
if pc = 24152 then
	inst <= x"02C0FFFF";
end if;
if pc = 24156 then
	inst <= x"82AC6420";
end if;
if pc = 24160 then
	inst <= x"02C00063";
end if;
if pc = 24164 then
	inst <= x"C47C0000";
end if;
if pc = 24168 then
	inst <= x"C45C0004";
end if;
if pc = 24172 then
	inst <= x"C43C0008";
end if;
if pc = 24176 then
	inst <= x"82AC6118";
end if;
if pc = 24180 then
	inst <= x"02C0030C";
end if;
if pc = 24184 then
	inst <= x"02E000C8";
end if;
if pc = 24188 then
	inst <= x"22AA0220";
end if;
if pc = 24192 then
	inst <= x"D0AEA000";
end if;
if pc = 24196 then
	inst <= x"C82C0000";
end if;
if pc = 24200 then
	inst <= x"C0EA0014";
end if;
if pc = 24204 then
	inst <= x"C84E0000";
end if;
if pc = 24208 then
	inst <= x"44224000";
end if;
if pc = 24212 then
	inst <= x"C84C0004";
end if;
if pc = 24216 then
	inst <= x"C0EA0014";
end if;
if pc = 24220 then
	inst <= x"C86E0004";
end if;
if pc = 24224 then
	inst <= x"44446000";
end if;
if pc = 24228 then
	inst <= x"C86C0008";
end if;
if pc = 24232 then
	inst <= x"C0CA0014";
end if;
if pc = 24236 then
	inst <= x"C88C0008";
end if;
if pc = 24240 then
	inst <= x"44668000";
end if;
if pc = 24244 then
	inst <= x"C0CA0004";
end if;
if pc = 24248 then
	inst <= x"02E00001";
end if;
if pc = 24252 then
	inst <= x"C49C000C";
end if;
if pc = 24256 then
	inst <= x"82CE5F14";
end if;
if pc = 24260 then
	inst <= x"02E00002";
end if;
if pc = 24264 then
	inst <= x"82CE5EF0";
end if;
if pc = 24268 then
	inst <= x"C17DFFFC";
end if;
if pc = 24272 then
	inst <= x"00460000";
end if;
if pc = 24276 then
	inst <= x"002A0000";
end if;
if pc = 24280 then
	inst <= x"03DC0018";
end if;
if pc = 24284 then
	inst <= x"037E000C";
end if;
if pc = 24288 then
	inst <= x"C57DFFFC";
end if;
if pc = 24292 then
	inst <= x"820034A0";
end if;
if pc = 24296 then
	inst <= x"07DC0018";
end if;
if pc = 24300 then
	inst <= x"82005F10";
end if;
if pc = 24304 then
	inst <= x"C17DFFFC";
end if;
if pc = 24308 then
	inst <= x"00460000";
end if;
if pc = 24312 then
	inst <= x"002A0000";
end if;
if pc = 24316 then
	inst <= x"03DC0018";
end if;
if pc = 24320 then
	inst <= x"037E000C";
end if;
if pc = 24324 then
	inst <= x"C57DFFFC";
end if;
if pc = 24328 then
	inst <= x"820032A4";
end if;
if pc = 24332 then
	inst <= x"07DC0018";
end if;
if pc = 24336 then
	inst <= x"82005FF4";
end if;
if pc = 24340 then
	inst <= x"02C00000";
end if;
if pc = 24344 then
	inst <= x"02E00001";
end if;
if pc = 24348 then
	inst <= x"03000002";
end if;
if pc = 24352 then
	inst <= x"CC3C0010";
end if;
if pc = 24356 then
	inst <= x"CC7C0018";
end if;
if pc = 24360 then
	inst <= x"CC5C0020";
end if;
if pc = 24364 then
	inst <= x"C4BC0028";
end if;
if pc = 24368 then
	inst <= x"C17DFFFC";
end if;
if pc = 24372 then
	inst <= x"008E0000";
end if;
if pc = 24376 then
	inst <= x"00460000";
end if;
if pc = 24380 then
	inst <= x"002A0000";
end if;
if pc = 24384 then
	inst <= x"00B00000";
end if;
if pc = 24388 then
	inst <= x"006C0000";
end if;
if pc = 24392 then
	inst <= x"03DC0034";
end if;
if pc = 24396 then
	inst <= x"037E000C";
end if;
if pc = 24400 then
	inst <= x"C57DFFFC";
end if;
if pc = 24404 then
	inst <= x"8200317C";
end if;
if pc = 24408 then
	inst <= x"07DC0034";
end if;
if pc = 24412 then
	inst <= x"82205F68";
end if;
if pc = 24416 then
	inst <= x"02200001";
end if;
if pc = 24420 then
	inst <= x"82005FF4";
end if;
if pc = 24424 then
	inst <= x"02600001";
end if;
if pc = 24428 then
	inst <= x"02800002";
end if;
if pc = 24432 then
	inst <= x"02A00000";
end if;
if pc = 24436 then
	inst <= x"C83C0020";
end if;
if pc = 24440 then
	inst <= x"C85C0018";
end if;
if pc = 24444 then
	inst <= x"C87C0010";
end if;
if pc = 24448 then
	inst <= x"C03C0028";
end if;
if pc = 24452 then
	inst <= x"C05C0000";
end if;
if pc = 24456 then
	inst <= x"C17DFFFC";
end if;
if pc = 24460 then
	inst <= x"03DC0034";
end if;
if pc = 24464 then
	inst <= x"037E000C";
end if;
if pc = 24468 then
	inst <= x"C57DFFFC";
end if;
if pc = 24472 then
	inst <= x"8200317C";
end if;
if pc = 24476 then
	inst <= x"07DC0034";
end if;
if pc = 24480 then
	inst <= x"82205FAC";
end if;
if pc = 24484 then
	inst <= x"02200002";
end if;
if pc = 24488 then
	inst <= x"82005FF4";
end if;
if pc = 24492 then
	inst <= x"02600002";
end if;
if pc = 24496 then
	inst <= x"02800000";
end if;
if pc = 24500 then
	inst <= x"02A00001";
end if;
if pc = 24504 then
	inst <= x"C83C0018";
end if;
if pc = 24508 then
	inst <= x"C85C0010";
end if;
if pc = 24512 then
	inst <= x"C87C0020";
end if;
if pc = 24516 then
	inst <= x"C03C0028";
end if;
if pc = 24520 then
	inst <= x"C05C0000";
end if;
if pc = 24524 then
	inst <= x"C17DFFFC";
end if;
if pc = 24528 then
	inst <= x"03DC0034";
end if;
if pc = 24532 then
	inst <= x"037E000C";
end if;
if pc = 24536 then
	inst <= x"C57DFFFC";
end if;
if pc = 24540 then
	inst <= x"8200317C";
end if;
if pc = 24544 then
	inst <= x"07DC0034";
end if;
if pc = 24548 then
	inst <= x"82205FF0";
end if;
if pc = 24552 then
	inst <= x"02200003";
end if;
if pc = 24556 then
	inst <= x"82005FF4";
end if;
if pc = 24560 then
	inst <= x"02200000";
end if;
if pc = 24564 then
	inst <= x"82206114";
end if;
if pc = 24568 then
	inst <= x"022002AC";
end if;
if pc = 24572 then
	inst <= x"C8220000";
end if;
if pc = 24576 then
	inst <= x"022002B4";
end if;
if pc = 24580 then
	inst <= x"C8420000";
end if;
if pc = 24584 then
	inst <= x"8E246010";
end if;
if pc = 24588 then
	inst <= x"82006110";
end if;
if pc = 24592 then
	inst <= x"C03C000C";
end if;
if pc = 24596 then
	inst <= x"C0420004";
end if;
if pc = 24600 then
	inst <= x"0260FFFF";
end if;
if pc = 24604 then
	inst <= x"82466110";
end if;
if pc = 24608 then
	inst <= x"026001E0";
end if;
if pc = 24612 then
	inst <= x"22440220";
end if;
if pc = 24616 then
	inst <= x"D0464000";
end if;
if pc = 24620 then
	inst <= x"02800000";
end if;
if pc = 24624 then
	inst <= x"C0BC0000";
end if;
if pc = 24628 then
	inst <= x"C47C002C";
end if;
if pc = 24632 then
	inst <= x"C17DFFFC";
end if;
if pc = 24636 then
	inst <= x"006A0000";
end if;
if pc = 24640 then
	inst <= x"00280000";
end if;
if pc = 24644 then
	inst <= x"03DC0038";
end if;
if pc = 24648 then
	inst <= x"037E000C";
end if;
if pc = 24652 then
	inst <= x"C57DFFFC";
end if;
if pc = 24656 then
	inst <= x"820057C8";
end if;
if pc = 24660 then
	inst <= x"07DC0038";
end if;
if pc = 24664 then
	inst <= x"C03C000C";
end if;
if pc = 24668 then
	inst <= x"C0420008";
end if;
if pc = 24672 then
	inst <= x"0260FFFF";
end if;
if pc = 24676 then
	inst <= x"8246610C";
end if;
if pc = 24680 then
	inst <= x"22440220";
end if;
if pc = 24684 then
	inst <= x"C07C002C";
end if;
if pc = 24688 then
	inst <= x"D0464000";
end if;
if pc = 24692 then
	inst <= x"02800000";
end if;
if pc = 24696 then
	inst <= x"C0BC0000";
end if;
if pc = 24700 then
	inst <= x"C17DFFFC";
end if;
if pc = 24704 then
	inst <= x"006A0000";
end if;
if pc = 24708 then
	inst <= x"00280000";
end if;
if pc = 24712 then
	inst <= x"03DC0038";
end if;
if pc = 24716 then
	inst <= x"037E000C";
end if;
if pc = 24720 then
	inst <= x"C57DFFFC";
end if;
if pc = 24724 then
	inst <= x"820057C8";
end if;
if pc = 24728 then
	inst <= x"07DC0038";
end if;
if pc = 24732 then
	inst <= x"C03C000C";
end if;
if pc = 24736 then
	inst <= x"C042000C";
end if;
if pc = 24740 then
	inst <= x"0260FFFF";
end if;
if pc = 24744 then
	inst <= x"82466108";
end if;
if pc = 24748 then
	inst <= x"22440220";
end if;
if pc = 24752 then
	inst <= x"C07C002C";
end if;
if pc = 24756 then
	inst <= x"D0464000";
end if;
if pc = 24760 then
	inst <= x"02600000";
end if;
if pc = 24764 then
	inst <= x"C09C0000";
end if;
if pc = 24768 then
	inst <= x"C17DFFFC";
end if;
if pc = 24772 then
	inst <= x"00260000";
end if;
if pc = 24776 then
	inst <= x"00680000";
end if;
if pc = 24780 then
	inst <= x"03DC0038";
end if;
if pc = 24784 then
	inst <= x"037E000C";
end if;
if pc = 24788 then
	inst <= x"C57DFFFC";
end if;
if pc = 24792 then
	inst <= x"820057C8";
end if;
if pc = 24796 then
	inst <= x"07DC0038";
end if;
if pc = 24800 then
	inst <= x"02200004";
end if;
if pc = 24804 then
	inst <= x"C05C000C";
end if;
if pc = 24808 then
	inst <= x"C07C0000";
end if;
if pc = 24812 then
	inst <= x"C17DFFFC";
end if;
if pc = 24816 then
	inst <= x"03DC0038";
end if;
if pc = 24820 then
	inst <= x"037E000C";
end if;
if pc = 24824 then
	inst <= x"C57DFFFC";
end if;
if pc = 24828 then
	inst <= x"82005CDC";
end if;
if pc = 24832 then
	inst <= x"07DC0038";
end if;
if pc = 24836 then
	inst <= x"82006108";
end if;
if pc = 24840 then
	inst <= x"8200610C";
end if;
if pc = 24844 then
	inst <= x"82006110";
end if;
if pc = 24848 then
	inst <= x"82006114";
end if;
if pc = 24852 then
	inst <= x"82006214";
end if;
if pc = 24856 then
	inst <= x"C0A80004";
end if;
if pc = 24860 then
	inst <= x"02C0FFFF";
end if;
if pc = 24864 then
	inst <= x"82AC6214";
end if;
if pc = 24868 then
	inst <= x"02C001E0";
end if;
if pc = 24872 then
	inst <= x"22AA0220";
end if;
if pc = 24876 then
	inst <= x"D0ACA000";
end if;
if pc = 24880 then
	inst <= x"02E00000";
end if;
if pc = 24884 then
	inst <= x"C4DC0030";
end if;
if pc = 24888 then
	inst <= x"C49C000C";
end if;
if pc = 24892 then
	inst <= x"C17DFFFC";
end if;
if pc = 24896 then
	inst <= x"004A0000";
end if;
if pc = 24900 then
	inst <= x"002E0000";
end if;
if pc = 24904 then
	inst <= x"03DC003C";
end if;
if pc = 24908 then
	inst <= x"037E000C";
end if;
if pc = 24912 then
	inst <= x"C57DFFFC";
end if;
if pc = 24916 then
	inst <= x"820057C8";
end if;
if pc = 24920 then
	inst <= x"07DC003C";
end if;
if pc = 24924 then
	inst <= x"C03C000C";
end if;
if pc = 24928 then
	inst <= x"C0420008";
end if;
if pc = 24932 then
	inst <= x"0260FFFF";
end if;
if pc = 24936 then
	inst <= x"82466210";
end if;
if pc = 24940 then
	inst <= x"22440220";
end if;
if pc = 24944 then
	inst <= x"C07C0030";
end if;
if pc = 24948 then
	inst <= x"D0464000";
end if;
if pc = 24952 then
	inst <= x"02800000";
end if;
if pc = 24956 then
	inst <= x"C0BC0000";
end if;
if pc = 24960 then
	inst <= x"C17DFFFC";
end if;
if pc = 24964 then
	inst <= x"006A0000";
end if;
if pc = 24968 then
	inst <= x"00280000";
end if;
if pc = 24972 then
	inst <= x"03DC003C";
end if;
if pc = 24976 then
	inst <= x"037E000C";
end if;
if pc = 24980 then
	inst <= x"C57DFFFC";
end if;
if pc = 24984 then
	inst <= x"820057C8";
end if;
if pc = 24988 then
	inst <= x"07DC003C";
end if;
if pc = 24992 then
	inst <= x"C03C000C";
end if;
if pc = 24996 then
	inst <= x"C042000C";
end if;
if pc = 25000 then
	inst <= x"0260FFFF";
end if;
if pc = 25004 then
	inst <= x"8246620C";
end if;
if pc = 25008 then
	inst <= x"22440220";
end if;
if pc = 25012 then
	inst <= x"C07C0030";
end if;
if pc = 25016 then
	inst <= x"D0464000";
end if;
if pc = 25020 then
	inst <= x"02600000";
end if;
if pc = 25024 then
	inst <= x"C09C0000";
end if;
if pc = 25028 then
	inst <= x"C17DFFFC";
end if;
if pc = 25032 then
	inst <= x"00260000";
end if;
if pc = 25036 then
	inst <= x"00680000";
end if;
if pc = 25040 then
	inst <= x"03DC003C";
end if;
if pc = 25044 then
	inst <= x"037E000C";
end if;
if pc = 25048 then
	inst <= x"C57DFFFC";
end if;
if pc = 25052 then
	inst <= x"820057C8";
end if;
if pc = 25056 then
	inst <= x"07DC003C";
end if;
if pc = 25060 then
	inst <= x"02200004";
end if;
if pc = 25064 then
	inst <= x"C05C000C";
end if;
if pc = 25068 then
	inst <= x"C07C0000";
end if;
if pc = 25072 then
	inst <= x"C17DFFFC";
end if;
if pc = 25076 then
	inst <= x"03DC003C";
end if;
if pc = 25080 then
	inst <= x"037E000C";
end if;
if pc = 25084 then
	inst <= x"C57DFFFC";
end if;
if pc = 25088 then
	inst <= x"82005CDC";
end if;
if pc = 25092 then
	inst <= x"07DC003C";
end if;
if pc = 25096 then
	inst <= x"8200620C";
end if;
if pc = 25100 then
	inst <= x"82006210";
end if;
if pc = 25104 then
	inst <= x"82006214";
end if;
if pc = 25108 then
	inst <= x"C03C0008";
end if;
if pc = 25112 then
	inst <= x"02220001";
end if;
if pc = 25116 then
	inst <= x"22420220";
end if;
if pc = 25120 then
	inst <= x"C07C0004";
end if;
if pc = 25124 then
	inst <= x"D0464000";
end if;
if pc = 25128 then
	inst <= x"C0840000";
end if;
if pc = 25132 then
	inst <= x"02A0FFFF";
end if;
if pc = 25136 then
	inst <= x"828A641C";
end if;
if pc = 25140 then
	inst <= x"02A00063";
end if;
if pc = 25144 then
	inst <= x"C43C0034";
end if;
if pc = 25148 then
	inst <= x"828A634C";
end if;
if pc = 25152 then
	inst <= x"02A0030C";
end if;
if pc = 25156 then
	inst <= x"C0DC0000";
end if;
if pc = 25160 then
	inst <= x"C45C0038";
end if;
if pc = 25164 then
	inst <= x"C17DFFFC";
end if;
if pc = 25168 then
	inst <= x"006A0000";
end if;
if pc = 25172 then
	inst <= x"004C0000";
end if;
if pc = 25176 then
	inst <= x"00280000";
end if;
if pc = 25180 then
	inst <= x"03DC0044";
end if;
if pc = 25184 then
	inst <= x"037E000C";
end if;
if pc = 25188 then
	inst <= x"C57DFFFC";
end if;
if pc = 25192 then
	inst <= x"820036D4";
end if;
if pc = 25196 then
	inst <= x"07DC0044";
end if;
if pc = 25200 then
	inst <= x"82206348";
end if;
if pc = 25204 then
	inst <= x"022002AC";
end if;
if pc = 25208 then
	inst <= x"C8220000";
end if;
if pc = 25212 then
	inst <= x"022002B4";
end if;
if pc = 25216 then
	inst <= x"C8420000";
end if;
if pc = 25220 then
	inst <= x"8E24628C";
end if;
if pc = 25224 then
	inst <= x"82006344";
end if;
if pc = 25228 then
	inst <= x"C03C0038";
end if;
if pc = 25232 then
	inst <= x"C0420004";
end if;
if pc = 25236 then
	inst <= x"0260FFFF";
end if;
if pc = 25240 then
	inst <= x"82466344";
end if;
if pc = 25244 then
	inst <= x"026001E0";
end if;
if pc = 25248 then
	inst <= x"22440220";
end if;
if pc = 25252 then
	inst <= x"D0464000";
end if;
if pc = 25256 then
	inst <= x"02800000";
end if;
if pc = 25260 then
	inst <= x"C0BC0000";
end if;
if pc = 25264 then
	inst <= x"C47C003C";
end if;
if pc = 25268 then
	inst <= x"C17DFFFC";
end if;
if pc = 25272 then
	inst <= x"006A0000";
end if;
if pc = 25276 then
	inst <= x"00280000";
end if;
if pc = 25280 then
	inst <= x"03DC0048";
end if;
if pc = 25284 then
	inst <= x"037E000C";
end if;
if pc = 25288 then
	inst <= x"C57DFFFC";
end if;
if pc = 25292 then
	inst <= x"820057C8";
end if;
if pc = 25296 then
	inst <= x"07DC0048";
end if;
if pc = 25300 then
	inst <= x"C03C0038";
end if;
if pc = 25304 then
	inst <= x"C0420008";
end if;
if pc = 25308 then
	inst <= x"0260FFFF";
end if;
if pc = 25312 then
	inst <= x"82466340";
end if;
if pc = 25316 then
	inst <= x"22440220";
end if;
if pc = 25320 then
	inst <= x"C07C003C";
end if;
if pc = 25324 then
	inst <= x"D0464000";
end if;
if pc = 25328 then
	inst <= x"02600000";
end if;
if pc = 25332 then
	inst <= x"C09C0000";
end if;
if pc = 25336 then
	inst <= x"C17DFFFC";
end if;
if pc = 25340 then
	inst <= x"00260000";
end if;
if pc = 25344 then
	inst <= x"00680000";
end if;
if pc = 25348 then
	inst <= x"03DC0048";
end if;
if pc = 25352 then
	inst <= x"037E000C";
end if;
if pc = 25356 then
	inst <= x"C57DFFFC";
end if;
if pc = 25360 then
	inst <= x"820057C8";
end if;
if pc = 25364 then
	inst <= x"07DC0048";
end if;
if pc = 25368 then
	inst <= x"02200003";
end if;
if pc = 25372 then
	inst <= x"C05C0038";
end if;
if pc = 25376 then
	inst <= x"C07C0000";
end if;
if pc = 25380 then
	inst <= x"C17DFFFC";
end if;
if pc = 25384 then
	inst <= x"03DC0048";
end if;
if pc = 25388 then
	inst <= x"037E000C";
end if;
if pc = 25392 then
	inst <= x"C57DFFFC";
end if;
if pc = 25396 then
	inst <= x"82005CDC";
end if;
if pc = 25400 then
	inst <= x"07DC0048";
end if;
if pc = 25404 then
	inst <= x"82006340";
end if;
if pc = 25408 then
	inst <= x"82006344";
end if;
if pc = 25412 then
	inst <= x"82006348";
end if;
if pc = 25416 then
	inst <= x"82006408";
end if;
if pc = 25420 then
	inst <= x"C0840004";
end if;
if pc = 25424 then
	inst <= x"02A0FFFF";
end if;
if pc = 25428 then
	inst <= x"828A6408";
end if;
if pc = 25432 then
	inst <= x"02A001E0";
end if;
if pc = 25436 then
	inst <= x"22880220";
end if;
if pc = 25440 then
	inst <= x"D08A8000";
end if;
if pc = 25444 then
	inst <= x"02C00000";
end if;
if pc = 25448 then
	inst <= x"C0FC0000";
end if;
if pc = 25452 then
	inst <= x"C4BC0040";
end if;
if pc = 25456 then
	inst <= x"C45C0038";
end if;
if pc = 25460 then
	inst <= x"C17DFFFC";
end if;
if pc = 25464 then
	inst <= x"006E0000";
end if;
if pc = 25468 then
	inst <= x"00480000";
end if;
if pc = 25472 then
	inst <= x"002C0000";
end if;
if pc = 25476 then
	inst <= x"03DC004C";
end if;
if pc = 25480 then
	inst <= x"037E000C";
end if;
if pc = 25484 then
	inst <= x"C57DFFFC";
end if;
if pc = 25488 then
	inst <= x"820057C8";
end if;
if pc = 25492 then
	inst <= x"07DC004C";
end if;
if pc = 25496 then
	inst <= x"C03C0038";
end if;
if pc = 25500 then
	inst <= x"C0420008";
end if;
if pc = 25504 then
	inst <= x"0260FFFF";
end if;
if pc = 25508 then
	inst <= x"82466404";
end if;
if pc = 25512 then
	inst <= x"22440220";
end if;
if pc = 25516 then
	inst <= x"C07C0040";
end if;
if pc = 25520 then
	inst <= x"D0464000";
end if;
if pc = 25524 then
	inst <= x"02600000";
end if;
if pc = 25528 then
	inst <= x"C09C0000";
end if;
if pc = 25532 then
	inst <= x"C17DFFFC";
end if;
if pc = 25536 then
	inst <= x"00260000";
end if;
if pc = 25540 then
	inst <= x"00680000";
end if;
if pc = 25544 then
	inst <= x"03DC004C";
end if;
if pc = 25548 then
	inst <= x"037E000C";
end if;
if pc = 25552 then
	inst <= x"C57DFFFC";
end if;
if pc = 25556 then
	inst <= x"820057C8";
end if;
if pc = 25560 then
	inst <= x"07DC004C";
end if;
if pc = 25564 then
	inst <= x"02200003";
end if;
if pc = 25568 then
	inst <= x"C05C0038";
end if;
if pc = 25572 then
	inst <= x"C07C0000";
end if;
if pc = 25576 then
	inst <= x"C17DFFFC";
end if;
if pc = 25580 then
	inst <= x"03DC004C";
end if;
if pc = 25584 then
	inst <= x"037E000C";
end if;
if pc = 25588 then
	inst <= x"C57DFFFC";
end if;
if pc = 25592 then
	inst <= x"82005CDC";
end if;
if pc = 25596 then
	inst <= x"07DC004C";
end if;
if pc = 25600 then
	inst <= x"82006404";
end if;
if pc = 25604 then
	inst <= x"82006408";
end if;
if pc = 25608 then
	inst <= x"C03C0034";
end if;
if pc = 25612 then
	inst <= x"02220001";
end if;
if pc = 25616 then
	inst <= x"C05C0004";
end if;
if pc = 25620 then
	inst <= x"C07C0000";
end if;
if pc = 25624 then
	inst <= x"82005E4C";
end if;
if pc = 25628 then
	inst <= x"C1FDFFFC";
end if;
if pc = 25632 then
	inst <= x"C1FDFFFC";
end if;
if pc = 25636 then
	inst <= x"C0860000";
end if;
if pc = 25640 then
	inst <= x"22A20220";
end if;
if pc = 25644 then
	inst <= x"D0A4A000";
end if;
if pc = 25648 then
	inst <= x"02C0FFFF";
end if;
if pc = 25652 then
	inst <= x"82AC6874";
end if;
if pc = 25656 then
	inst <= x"02C000C8";
end if;
if pc = 25660 then
	inst <= x"22EA0220";
end if;
if pc = 25664 then
	inst <= x"D0ECE000";
end if;
if pc = 25668 then
	inst <= x"C10E0028";
end if;
if pc = 25672 then
	inst <= x"C8300000";
end if;
if pc = 25676 then
	inst <= x"C8500004";
end if;
if pc = 25680 then
	inst <= x"C8700008";
end if;
if pc = 25684 then
	inst <= x"C1260004";
end if;
if pc = 25688 then
	inst <= x"234A0220";
end if;
if pc = 25692 then
	inst <= x"D1334000";
end if;
if pc = 25696 then
	inst <= x"C14E0004";
end if;
if pc = 25700 then
	inst <= x"C49C0000";
end if;
if pc = 25704 then
	inst <= x"02800001";
end if;
if pc = 25708 then
	inst <= x"C47C0004";
end if;
if pc = 25712 then
	inst <= x"C45C0008";
end if;
if pc = 25716 then
	inst <= x"C43C000C";
end if;
if pc = 25720 then
	inst <= x"C4DC0010";
end if;
if pc = 25724 then
	inst <= x"C4BC0014";
end if;
if pc = 25728 then
	inst <= x"834864E0";
end if;
if pc = 25732 then
	inst <= x"02800002";
end if;
if pc = 25736 then
	inst <= x"834864B4";
end if;
if pc = 25740 then
	inst <= x"C17DFFFC";
end if;
if pc = 25744 then
	inst <= x"00700000";
end if;
if pc = 25748 then
	inst <= x"00520000";
end if;
if pc = 25752 then
	inst <= x"002E0000";
end if;
if pc = 25756 then
	inst <= x"03DC0020";
end if;
if pc = 25760 then
	inst <= x"037E000C";
end if;
if pc = 25764 then
	inst <= x"C57DFFFC";
end if;
if pc = 25768 then
	inst <= x"82003BD4";
end if;
if pc = 25772 then
	inst <= x"07DC0020";
end if;
if pc = 25776 then
	inst <= x"820064DC";
end if;
if pc = 25780 then
	inst <= x"C8320000";
end if;
if pc = 25784 then
	inst <= x"8E2064C4";
end if;
if pc = 25788 then
	inst <= x"02200000";
end if;
if pc = 25792 then
	inst <= x"820064DC";
end if;
if pc = 25796 then
	inst <= x"028002AC";
end if;
if pc = 25800 then
	inst <= x"C8320000";
end if;
if pc = 25804 then
	inst <= x"C850000C";
end if;
if pc = 25808 then
	inst <= x"48224000";
end if;
if pc = 25812 then
	inst <= x"CC280000";
end if;
if pc = 25816 then
	inst <= x"02200001";
end if;
if pc = 25820 then
	inst <= x"82006508";
end if;
if pc = 25824 then
	inst <= x"C0860000";
end if;
if pc = 25828 then
	inst <= x"C17DFFFC";
end if;
if pc = 25832 then
	inst <= x"00720000";
end if;
if pc = 25836 then
	inst <= x"00480000";
end if;
if pc = 25840 then
	inst <= x"002E0000";
end if;
if pc = 25844 then
	inst <= x"03DC0020";
end if;
if pc = 25848 then
	inst <= x"037E000C";
end if;
if pc = 25852 then
	inst <= x"C57DFFFC";
end if;
if pc = 25856 then
	inst <= x"8200389C";
end if;
if pc = 25860 then
	inst <= x"07DC0020";
end if;
if pc = 25864 then
	inst <= x"82206844";
end if;
if pc = 25868 then
	inst <= x"024002AC";
end if;
if pc = 25872 then
	inst <= x"C8240000";
end if;
if pc = 25876 then
	inst <= x"8E02651C";
end if;
if pc = 25880 then
	inst <= x"82006830";
end if;
if pc = 25884 then
	inst <= x"024002B4";
end if;
if pc = 25888 then
	inst <= x"C8440000";
end if;
if pc = 25892 then
	inst <= x"8E24652C";
end if;
if pc = 25896 then
	inst <= x"82006830";
end if;
if pc = 25900 then
	inst <= x"C8400074";
end if;
if pc = 25904 then
	inst <= x"40224000";
end if;
if pc = 25908 then
	inst <= x"C07C0000";
end if;
if pc = 25912 then
	inst <= x"C8460000";
end if;
if pc = 25916 then
	inst <= x"48442000";
end if;
if pc = 25920 then
	inst <= x"02800318";
end if;
if pc = 25924 then
	inst <= x"C8680000";
end if;
if pc = 25928 then
	inst <= x"40446000";
end if;
if pc = 25932 then
	inst <= x"C8660004";
end if;
if pc = 25936 then
	inst <= x"48662000";
end if;
if pc = 25940 then
	inst <= x"C8880004";
end if;
if pc = 25944 then
	inst <= x"40668000";
end if;
if pc = 25948 then
	inst <= x"C8860008";
end if;
if pc = 25952 then
	inst <= x"48882000";
end if;
if pc = 25956 then
	inst <= x"C8A80008";
end if;
if pc = 25960 then
	inst <= x"4088A000";
end if;
if pc = 25964 then
	inst <= x"C07C0008";
end if;
if pc = 25968 then
	inst <= x"C0860000";
end if;
if pc = 25972 then
	inst <= x"02A0FFFF";
end if;
if pc = 25976 then
	inst <= x"C43C0018";
end if;
if pc = 25980 then
	inst <= x"CC9C0020";
end if;
if pc = 25984 then
	inst <= x"CC7C0028";
end if;
if pc = 25988 then
	inst <= x"CC5C0030";
end if;
if pc = 25992 then
	inst <= x"C45C0038";
end if;
if pc = 25996 then
	inst <= x"CC3C0040";
end if;
if pc = 26000 then
	inst <= x"828A67E4";
end if;
if pc = 26004 then
	inst <= x"22880220";
end if;
if pc = 26008 then
	inst <= x"C0BC0010";
end if;
if pc = 26012 then
	inst <= x"D08A8000";
end if;
if pc = 26016 then
	inst <= x"C17DFFFC";
end if;
if pc = 26020 then
	inst <= x"00280000";
end if;
if pc = 26024 then
	inst <= x"40204000";
end if;
if pc = 26028 then
	inst <= x"40406000";
end if;
if pc = 26032 then
	inst <= x"40608000";
end if;
if pc = 26036 then
	inst <= x"03DC0050";
end if;
if pc = 26040 then
	inst <= x"037E000C";
end if;
if pc = 26044 then
	inst <= x"C57DFFFC";
end if;
if pc = 26048 then
	inst <= x"82004860";
end if;
if pc = 26052 then
	inst <= x"07DC0050";
end if;
if pc = 26056 then
	inst <= x"822065D4";
end if;
if pc = 26060 then
	inst <= x"02200000";
end if;
if pc = 26064 then
	inst <= x"820067E0";
end if;
if pc = 26068 then
	inst <= x"C05C0008";
end if;
if pc = 26072 then
	inst <= x"C0240004";
end if;
if pc = 26076 then
	inst <= x"0260FFFF";
end if;
if pc = 26080 then
	inst <= x"822667DC";
end if;
if pc = 26084 then
	inst <= x"22220220";
end if;
if pc = 26088 then
	inst <= x"C07C0010";
end if;
if pc = 26092 then
	inst <= x"D0262000";
end if;
if pc = 26096 then
	inst <= x"C0820014";
end if;
if pc = 26100 then
	inst <= x"C8280000";
end if;
if pc = 26104 then
	inst <= x"C85C0030";
end if;
if pc = 26108 then
	inst <= x"44242000";
end if;
if pc = 26112 then
	inst <= x"C0820014";
end if;
if pc = 26116 then
	inst <= x"C8680004";
end if;
if pc = 26120 then
	inst <= x"C89C0028";
end if;
if pc = 26124 then
	inst <= x"44686000";
end if;
if pc = 26128 then
	inst <= x"C0820014";
end if;
if pc = 26132 then
	inst <= x"C8A80008";
end if;
if pc = 26136 then
	inst <= x"C8DC0020";
end if;
if pc = 26140 then
	inst <= x"44ACA000";
end if;
if pc = 26144 then
	inst <= x"C0820004";
end if;
if pc = 26148 then
	inst <= x"02A00001";
end if;
if pc = 26152 then
	inst <= x"828A66C0";
end if;
if pc = 26156 then
	inst <= x"02A00002";
end if;
if pc = 26160 then
	inst <= x"828A6658";
end if;
if pc = 26164 then
	inst <= x"C17DFFFC";
end if;
if pc = 26168 then
	inst <= x"40406000";
end if;
if pc = 26172 then
	inst <= x"4060A000";
end if;
if pc = 26176 then
	inst <= x"03DC0050";
end if;
if pc = 26180 then
	inst <= x"037E000C";
end if;
if pc = 26184 then
	inst <= x"C57DFFFC";
end if;
if pc = 26188 then
	inst <= x"82004780";
end if;
if pc = 26192 then
	inst <= x"07DC0050";
end if;
if pc = 26196 then
	inst <= x"820066BC";
end if;
if pc = 26200 then
	inst <= x"C0820010";
end if;
if pc = 26204 then
	inst <= x"C8E80000";
end if;
if pc = 26208 then
	inst <= x"482E2000";
end if;
if pc = 26212 then
	inst <= x"C8E80004";
end if;
if pc = 26216 then
	inst <= x"486E6000";
end if;
if pc = 26220 then
	inst <= x"40226000";
end if;
if pc = 26224 then
	inst <= x"C8680008";
end if;
if pc = 26228 then
	inst <= x"4866A000";
end if;
if pc = 26232 then
	inst <= x"40226000";
end if;
if pc = 26236 then
	inst <= x"C0220018";
end if;
if pc = 26240 then
	inst <= x"8E20668C";
end if;
if pc = 26244 then
	inst <= x"02800000";
end if;
if pc = 26248 then
	inst <= x"82006690";
end if;
if pc = 26252 then
	inst <= x"02800001";
end if;
if pc = 26256 then
	inst <= x"822066A8";
end if;
if pc = 26260 then
	inst <= x"8E2066A0";
end if;
if pc = 26264 then
	inst <= x"02200001";
end if;
if pc = 26268 then
	inst <= x"820066A4";
end if;
if pc = 26272 then
	inst <= x"02200000";
end if;
if pc = 26276 then
	inst <= x"820066AC";
end if;
if pc = 26280 then
	inst <= x"00280000";
end if;
if pc = 26284 then
	inst <= x"822066B8";
end if;
if pc = 26288 then
	inst <= x"02200000";
end if;
if pc = 26292 then
	inst <= x"820066BC";
end if;
if pc = 26296 then
	inst <= x"02200001";
end if;
if pc = 26300 then
	inst <= x"8200674C";
end if;
if pc = 26304 then
	inst <= x"8E2066C8";
end if;
if pc = 26308 then
	inst <= x"820066CC";
end if;
if pc = 26312 then
	inst <= x"44202000";
end if;
if pc = 26316 then
	inst <= x"C0820010";
end if;
if pc = 26320 then
	inst <= x"C8E80000";
end if;
if pc = 26324 then
	inst <= x"8E2E66E0";
end if;
if pc = 26328 then
	inst <= x"02800000";
end if;
if pc = 26332 then
	inst <= x"8200672C";
end if;
if pc = 26336 then
	inst <= x"8E6066EC";
end if;
if pc = 26340 then
	inst <= x"40206000";
end if;
if pc = 26344 then
	inst <= x"820066F0";
end if;
if pc = 26348 then
	inst <= x"44206000";
end if;
if pc = 26352 then
	inst <= x"C0820010";
end if;
if pc = 26356 then
	inst <= x"C8680004";
end if;
if pc = 26360 then
	inst <= x"8E266704";
end if;
if pc = 26364 then
	inst <= x"02800000";
end if;
if pc = 26368 then
	inst <= x"8200672C";
end if;
if pc = 26372 then
	inst <= x"8EA06710";
end if;
if pc = 26376 then
	inst <= x"4020A000";
end if;
if pc = 26380 then
	inst <= x"82006714";
end if;
if pc = 26384 then
	inst <= x"4420A000";
end if;
if pc = 26388 then
	inst <= x"C0820010";
end if;
if pc = 26392 then
	inst <= x"C8680008";
end if;
if pc = 26396 then
	inst <= x"8E266728";
end if;
if pc = 26400 then
	inst <= x"02800000";
end if;
if pc = 26404 then
	inst <= x"8200672C";
end if;
if pc = 26408 then
	inst <= x"02800001";
end if;
if pc = 26412 then
	inst <= x"82806738";
end if;
if pc = 26416 then
	inst <= x"C0220018";
end if;
if pc = 26420 then
	inst <= x"8200674C";
end if;
if pc = 26424 then
	inst <= x"C0220018";
end if;
if pc = 26428 then
	inst <= x"82206748";
end if;
if pc = 26432 then
	inst <= x"02200000";
end if;
if pc = 26436 then
	inst <= x"8200674C";
end if;
if pc = 26440 then
	inst <= x"02200001";
end if;
if pc = 26444 then
	inst <= x"82206758";
end if;
if pc = 26448 then
	inst <= x"02200000";
end if;
if pc = 26452 then
	inst <= x"820067D8";
end if;
if pc = 26456 then
	inst <= x"C05C0008";
end if;
if pc = 26460 then
	inst <= x"C0240008";
end if;
if pc = 26464 then
	inst <= x"0260FFFF";
end if;
if pc = 26468 then
	inst <= x"822667D4";
end if;
if pc = 26472 then
	inst <= x"22220220";
end if;
if pc = 26476 then
	inst <= x"C07C0010";
end if;
if pc = 26480 then
	inst <= x"D0262000";
end if;
if pc = 26484 then
	inst <= x"C83C0030";
end if;
if pc = 26488 then
	inst <= x"C85C0028";
end if;
if pc = 26492 then
	inst <= x"C87C0020";
end if;
if pc = 26496 then
	inst <= x"C17DFFFC";
end if;
if pc = 26500 then
	inst <= x"03DC0050";
end if;
if pc = 26504 then
	inst <= x"037E000C";
end if;
if pc = 26508 then
	inst <= x"C57DFFFC";
end if;
if pc = 26512 then
	inst <= x"82004860";
end if;
if pc = 26516 then
	inst <= x"07DC0050";
end if;
if pc = 26520 then
	inst <= x"822067A4";
end if;
if pc = 26524 then
	inst <= x"02200000";
end if;
if pc = 26528 then
	inst <= x"820067D0";
end if;
if pc = 26532 then
	inst <= x"02200003";
end if;
if pc = 26536 then
	inst <= x"C83C0030";
end if;
if pc = 26540 then
	inst <= x"C85C0028";
end if;
if pc = 26544 then
	inst <= x"C87C0020";
end if;
if pc = 26548 then
	inst <= x"C05C0008";
end if;
if pc = 26552 then
	inst <= x"C17DFFFC";
end if;
if pc = 26556 then
	inst <= x"03DC0050";
end if;
if pc = 26560 then
	inst <= x"037E000C";
end if;
if pc = 26564 then
	inst <= x"C57DFFFC";
end if;
if pc = 26568 then
	inst <= x"82004A0C";
end if;
if pc = 26572 then
	inst <= x"07DC0050";
end if;
if pc = 26576 then
	inst <= x"820067D8";
end if;
if pc = 26580 then
	inst <= x"02200001";
end if;
if pc = 26584 then
	inst <= x"820067E0";
end if;
if pc = 26588 then
	inst <= x"02200001";
end if;
if pc = 26592 then
	inst <= x"820067E8";
end if;
if pc = 26596 then
	inst <= x"02200001";
end if;
if pc = 26600 then
	inst <= x"82206830";
end if;
if pc = 26604 then
	inst <= x"C03C0038";
end if;
if pc = 26608 then
	inst <= x"C83C0040";
end if;
if pc = 26612 then
	inst <= x"CC220000";
end if;
if pc = 26616 then
	inst <= x"022002B8";
end if;
if pc = 26620 then
	inst <= x"C83C0030";
end if;
if pc = 26624 then
	inst <= x"CC220000";
end if;
if pc = 26628 then
	inst <= x"C83C0028";
end if;
if pc = 26632 then
	inst <= x"CC220004";
end if;
if pc = 26636 then
	inst <= x"C83C0020";
end if;
if pc = 26640 then
	inst <= x"CC220008";
end if;
if pc = 26644 then
	inst <= x"022002C4";
end if;
if pc = 26648 then
	inst <= x"C05C0014";
end if;
if pc = 26652 then
	inst <= x"C4420000";
end if;
if pc = 26656 then
	inst <= x"022002B0";
end if;
if pc = 26660 then
	inst <= x"C05C0018";
end if;
if pc = 26664 then
	inst <= x"C4420000";
end if;
if pc = 26668 then
	inst <= x"82006830";
end if;
if pc = 26672 then
	inst <= x"C03C000C";
end if;
if pc = 26676 then
	inst <= x"02220001";
end if;
if pc = 26680 then
	inst <= x"C05C0008";
end if;
if pc = 26684 then
	inst <= x"C07C0004";
end if;
if pc = 26688 then
	inst <= x"82006424";
end if;
if pc = 26692 then
	inst <= x"C03C0014";
end if;
if pc = 26696 then
	inst <= x"22220220";
end if;
if pc = 26700 then
	inst <= x"C05C0010";
end if;
if pc = 26704 then
	inst <= x"D0242000";
end if;
if pc = 26708 then
	inst <= x"C0220018";
end if;
if pc = 26712 then
	inst <= x"82206870";
end if;
if pc = 26716 then
	inst <= x"C03C000C";
end if;
if pc = 26720 then
	inst <= x"02220001";
end if;
if pc = 26724 then
	inst <= x"C05C0008";
end if;
if pc = 26728 then
	inst <= x"C07C0004";
end if;
if pc = 26732 then
	inst <= x"82006424";
end if;
if pc = 26736 then
	inst <= x"C1FDFFFC";
end if;
if pc = 26740 then
	inst <= x"C1FDFFFC";
end if;
if pc = 26744 then
	inst <= x"22820220";
end if;
if pc = 26748 then
	inst <= x"D0848000";
end if;
if pc = 26752 then
	inst <= x"02A0FFFF";
end if;
if pc = 26756 then
	inst <= x"828A69E4";
end if;
if pc = 26760 then
	inst <= x"02A001E0";
end if;
if pc = 26764 then
	inst <= x"22880220";
end if;
if pc = 26768 then
	inst <= x"D08A8000";
end if;
if pc = 26772 then
	inst <= x"02C00000";
end if;
if pc = 26776 then
	inst <= x"C47C0000";
end if;
if pc = 26780 then
	inst <= x"C4BC0004";
end if;
if pc = 26784 then
	inst <= x"C45C0008";
end if;
if pc = 26788 then
	inst <= x"C43C000C";
end if;
if pc = 26792 then
	inst <= x"C17DFFFC";
end if;
if pc = 26796 then
	inst <= x"00480000";
end if;
if pc = 26800 then
	inst <= x"002C0000";
end if;
if pc = 26804 then
	inst <= x"03DC0018";
end if;
if pc = 26808 then
	inst <= x"037E000C";
end if;
if pc = 26812 then
	inst <= x"C57DFFFC";
end if;
if pc = 26816 then
	inst <= x"82006424";
end if;
if pc = 26820 then
	inst <= x"07DC0018";
end if;
if pc = 26824 then
	inst <= x"C03C000C";
end if;
if pc = 26828 then
	inst <= x"02220001";
end if;
if pc = 26832 then
	inst <= x"22420220";
end if;
if pc = 26836 then
	inst <= x"C07C0008";
end if;
if pc = 26840 then
	inst <= x"D0464000";
end if;
if pc = 26844 then
	inst <= x"0280FFFF";
end if;
if pc = 26848 then
	inst <= x"824869E0";
end if;
if pc = 26852 then
	inst <= x"22440220";
end if;
if pc = 26856 then
	inst <= x"C09C0004";
end if;
if pc = 26860 then
	inst <= x"D0484000";
end if;
if pc = 26864 then
	inst <= x"02A00000";
end if;
if pc = 26868 then
	inst <= x"C0DC0000";
end if;
if pc = 26872 then
	inst <= x"C43C0010";
end if;
if pc = 26876 then
	inst <= x"C17DFFFC";
end if;
if pc = 26880 then
	inst <= x"006C0000";
end if;
if pc = 26884 then
	inst <= x"002A0000";
end if;
if pc = 26888 then
	inst <= x"03DC001C";
end if;
if pc = 26892 then
	inst <= x"037E000C";
end if;
if pc = 26896 then
	inst <= x"C57DFFFC";
end if;
if pc = 26900 then
	inst <= x"82006424";
end if;
if pc = 26904 then
	inst <= x"07DC001C";
end if;
if pc = 26908 then
	inst <= x"C03C0010";
end if;
if pc = 26912 then
	inst <= x"02220001";
end if;
if pc = 26916 then
	inst <= x"22420220";
end if;
if pc = 26920 then
	inst <= x"C07C0008";
end if;
if pc = 26924 then
	inst <= x"D0464000";
end if;
if pc = 26928 then
	inst <= x"0280FFFF";
end if;
if pc = 26932 then
	inst <= x"824869DC";
end if;
if pc = 26936 then
	inst <= x"22440220";
end if;
if pc = 26940 then
	inst <= x"C09C0004";
end if;
if pc = 26944 then
	inst <= x"D0484000";
end if;
if pc = 26948 then
	inst <= x"02A00000";
end if;
if pc = 26952 then
	inst <= x"C0DC0000";
end if;
if pc = 26956 then
	inst <= x"C43C0014";
end if;
if pc = 26960 then
	inst <= x"C17DFFFC";
end if;
if pc = 26964 then
	inst <= x"006C0000";
end if;
if pc = 26968 then
	inst <= x"002A0000";
end if;
if pc = 26972 then
	inst <= x"03DC0020";
end if;
if pc = 26976 then
	inst <= x"037E000C";
end if;
if pc = 26980 then
	inst <= x"C57DFFFC";
end if;
if pc = 26984 then
	inst <= x"82006424";
end if;
if pc = 26988 then
	inst <= x"07DC0020";
end if;
if pc = 26992 then
	inst <= x"C03C0014";
end if;
if pc = 26996 then
	inst <= x"02220001";
end if;
if pc = 27000 then
	inst <= x"22420220";
end if;
if pc = 27004 then
	inst <= x"C07C0008";
end if;
if pc = 27008 then
	inst <= x"D0464000";
end if;
if pc = 27012 then
	inst <= x"0280FFFF";
end if;
if pc = 27016 then
	inst <= x"824869D8";
end if;
if pc = 27020 then
	inst <= x"22440220";
end if;
if pc = 27024 then
	inst <= x"C09C0004";
end if;
if pc = 27028 then
	inst <= x"D0484000";
end if;
if pc = 27032 then
	inst <= x"02800000";
end if;
if pc = 27036 then
	inst <= x"C0BC0000";
end if;
if pc = 27040 then
	inst <= x"C43C0018";
end if;
if pc = 27044 then
	inst <= x"C17DFFFC";
end if;
if pc = 27048 then
	inst <= x"006A0000";
end if;
if pc = 27052 then
	inst <= x"00280000";
end if;
if pc = 27056 then
	inst <= x"03DC0024";
end if;
if pc = 27060 then
	inst <= x"037E000C";
end if;
if pc = 27064 then
	inst <= x"C57DFFFC";
end if;
if pc = 27068 then
	inst <= x"82006424";
end if;
if pc = 27072 then
	inst <= x"07DC0024";
end if;
if pc = 27076 then
	inst <= x"C03C0018";
end if;
if pc = 27080 then
	inst <= x"02220001";
end if;
if pc = 27084 then
	inst <= x"C05C0008";
end if;
if pc = 27088 then
	inst <= x"C07C0000";
end if;
if pc = 27092 then
	inst <= x"82006878";
end if;
if pc = 27096 then
	inst <= x"C1FDFFFC";
end if;
if pc = 27100 then
	inst <= x"C1FDFFFC";
end if;
if pc = 27104 then
	inst <= x"C1FDFFFC";
end if;
if pc = 27108 then
	inst <= x"C1FDFFFC";
end if;
if pc = 27112 then
	inst <= x"22820220";
end if;
if pc = 27116 then
	inst <= x"D0848000";
end if;
if pc = 27120 then
	inst <= x"C0A80000";
end if;
if pc = 27124 then
	inst <= x"02C0FFFF";
end if;
if pc = 27128 then
	inst <= x"82AC6F88";
end if;
if pc = 27132 then
	inst <= x"02C00063";
end if;
if pc = 27136 then
	inst <= x"C47C0000";
end if;
if pc = 27140 then
	inst <= x"C45C0004";
end if;
if pc = 27144 then
	inst <= x"C43C0008";
end if;
if pc = 27148 then
	inst <= x"82AC6BF0";
end if;
if pc = 27152 then
	inst <= x"02C000C8";
end if;
if pc = 27156 then
	inst <= x"22EA0220";
end if;
if pc = 27160 then
	inst <= x"D0CCE000";
end if;
if pc = 27164 then
	inst <= x"C0EC0028";
end if;
if pc = 27168 then
	inst <= x"C82E0000";
end if;
if pc = 27172 then
	inst <= x"C84E0004";
end if;
if pc = 27176 then
	inst <= x"C86E0008";
end if;
if pc = 27180 then
	inst <= x"C1060004";
end if;
if pc = 27184 then
	inst <= x"22AA0220";
end if;
if pc = 27188 then
	inst <= x"D0B0A000";
end if;
if pc = 27192 then
	inst <= x"C10C0004";
end if;
if pc = 27196 then
	inst <= x"03200001";
end if;
if pc = 27200 then
	inst <= x"C49C000C";
end if;
if pc = 27204 then
	inst <= x"83126AA4";
end if;
if pc = 27208 then
	inst <= x"03200002";
end if;
if pc = 27212 then
	inst <= x"83126A78";
end if;
if pc = 27216 then
	inst <= x"C17DFFFC";
end if;
if pc = 27220 then
	inst <= x"006E0000";
end if;
if pc = 27224 then
	inst <= x"004A0000";
end if;
if pc = 27228 then
	inst <= x"002C0000";
end if;
if pc = 27232 then
	inst <= x"03DC0018";
end if;
if pc = 27236 then
	inst <= x"037E000C";
end if;
if pc = 27240 then
	inst <= x"C57DFFFC";
end if;
if pc = 27244 then
	inst <= x"82003BD4";
end if;
if pc = 27248 then
	inst <= x"07DC0018";
end if;
if pc = 27252 then
	inst <= x"82006AA0";
end if;
if pc = 27256 then
	inst <= x"C82A0000";
end if;
if pc = 27260 then
	inst <= x"8E206A88";
end if;
if pc = 27264 then
	inst <= x"02200000";
end if;
if pc = 27268 then
	inst <= x"82006AA0";
end if;
if pc = 27272 then
	inst <= x"02C002AC";
end if;
if pc = 27276 then
	inst <= x"C82A0000";
end if;
if pc = 27280 then
	inst <= x"C84E000C";
end if;
if pc = 27284 then
	inst <= x"48224000";
end if;
if pc = 27288 then
	inst <= x"CC2C0000";
end if;
if pc = 27292 then
	inst <= x"02200001";
end if;
if pc = 27296 then
	inst <= x"82006ACC";
end if;
if pc = 27300 then
	inst <= x"C0E60000";
end if;
if pc = 27304 then
	inst <= x"C17DFFFC";
end if;
if pc = 27308 then
	inst <= x"006A0000";
end if;
if pc = 27312 then
	inst <= x"004E0000";
end if;
if pc = 27316 then
	inst <= x"002C0000";
end if;
if pc = 27320 then
	inst <= x"03DC0018";
end if;
if pc = 27324 then
	inst <= x"037E000C";
end if;
if pc = 27328 then
	inst <= x"C57DFFFC";
end if;
if pc = 27332 then
	inst <= x"8200389C";
end if;
if pc = 27336 then
	inst <= x"07DC0018";
end if;
if pc = 27340 then
	inst <= x"82206BEC";
end if;
if pc = 27344 then
	inst <= x"022002AC";
end if;
if pc = 27348 then
	inst <= x"C8220000";
end if;
if pc = 27352 then
	inst <= x"022002B4";
end if;
if pc = 27356 then
	inst <= x"C8420000";
end if;
if pc = 27360 then
	inst <= x"8E246AE8";
end if;
if pc = 27364 then
	inst <= x"82006BE8";
end if;
if pc = 27368 then
	inst <= x"C03C000C";
end if;
if pc = 27372 then
	inst <= x"C0420004";
end if;
if pc = 27376 then
	inst <= x"0260FFFF";
end if;
if pc = 27380 then
	inst <= x"82466BE8";
end if;
if pc = 27384 then
	inst <= x"026001E0";
end if;
if pc = 27388 then
	inst <= x"22440220";
end if;
if pc = 27392 then
	inst <= x"D0464000";
end if;
if pc = 27396 then
	inst <= x"02800000";
end if;
if pc = 27400 then
	inst <= x"C0BC0000";
end if;
if pc = 27404 then
	inst <= x"C47C0010";
end if;
if pc = 27408 then
	inst <= x"C17DFFFC";
end if;
if pc = 27412 then
	inst <= x"006A0000";
end if;
if pc = 27416 then
	inst <= x"00280000";
end if;
if pc = 27420 then
	inst <= x"03DC001C";
end if;
if pc = 27424 then
	inst <= x"037E000C";
end if;
if pc = 27428 then
	inst <= x"C57DFFFC";
end if;
if pc = 27432 then
	inst <= x"82006424";
end if;
if pc = 27436 then
	inst <= x"07DC001C";
end if;
if pc = 27440 then
	inst <= x"C03C000C";
end if;
if pc = 27444 then
	inst <= x"C0420008";
end if;
if pc = 27448 then
	inst <= x"0260FFFF";
end if;
if pc = 27452 then
	inst <= x"82466BE4";
end if;
if pc = 27456 then
	inst <= x"22440220";
end if;
if pc = 27460 then
	inst <= x"C07C0010";
end if;
if pc = 27464 then
	inst <= x"D0464000";
end if;
if pc = 27468 then
	inst <= x"02800000";
end if;
if pc = 27472 then
	inst <= x"C0BC0000";
end if;
if pc = 27476 then
	inst <= x"C17DFFFC";
end if;
if pc = 27480 then
	inst <= x"006A0000";
end if;
if pc = 27484 then
	inst <= x"00280000";
end if;
if pc = 27488 then
	inst <= x"03DC001C";
end if;
if pc = 27492 then
	inst <= x"037E000C";
end if;
if pc = 27496 then
	inst <= x"C57DFFFC";
end if;
if pc = 27500 then
	inst <= x"82006424";
end if;
if pc = 27504 then
	inst <= x"07DC001C";
end if;
if pc = 27508 then
	inst <= x"C03C000C";
end if;
if pc = 27512 then
	inst <= x"C042000C";
end if;
if pc = 27516 then
	inst <= x"0260FFFF";
end if;
if pc = 27520 then
	inst <= x"82466BE0";
end if;
if pc = 27524 then
	inst <= x"22440220";
end if;
if pc = 27528 then
	inst <= x"C07C0010";
end if;
if pc = 27532 then
	inst <= x"D0464000";
end if;
if pc = 27536 then
	inst <= x"02600000";
end if;
if pc = 27540 then
	inst <= x"C09C0000";
end if;
if pc = 27544 then
	inst <= x"C17DFFFC";
end if;
if pc = 27548 then
	inst <= x"00260000";
end if;
if pc = 27552 then
	inst <= x"00680000";
end if;
if pc = 27556 then
	inst <= x"03DC001C";
end if;
if pc = 27560 then
	inst <= x"037E000C";
end if;
if pc = 27564 then
	inst <= x"C57DFFFC";
end if;
if pc = 27568 then
	inst <= x"82006424";
end if;
if pc = 27572 then
	inst <= x"07DC001C";
end if;
if pc = 27576 then
	inst <= x"02200004";
end if;
if pc = 27580 then
	inst <= x"C05C000C";
end if;
if pc = 27584 then
	inst <= x"C07C0000";
end if;
if pc = 27588 then
	inst <= x"C17DFFFC";
end if;
if pc = 27592 then
	inst <= x"03DC001C";
end if;
if pc = 27596 then
	inst <= x"037E000C";
end if;
if pc = 27600 then
	inst <= x"C57DFFFC";
end if;
if pc = 27604 then
	inst <= x"82006878";
end if;
if pc = 27608 then
	inst <= x"07DC001C";
end if;
if pc = 27612 then
	inst <= x"82006BE0";
end if;
if pc = 27616 then
	inst <= x"82006BE4";
end if;
if pc = 27620 then
	inst <= x"82006BE8";
end if;
if pc = 27624 then
	inst <= x"82006BEC";
end if;
if pc = 27628 then
	inst <= x"82006CEC";
end if;
if pc = 27632 then
	inst <= x"C0A80004";
end if;
if pc = 27636 then
	inst <= x"02C0FFFF";
end if;
if pc = 27640 then
	inst <= x"82AC6CEC";
end if;
if pc = 27644 then
	inst <= x"02C001E0";
end if;
if pc = 27648 then
	inst <= x"22AA0220";
end if;
if pc = 27652 then
	inst <= x"D0ACA000";
end if;
if pc = 27656 then
	inst <= x"02E00000";
end if;
if pc = 27660 then
	inst <= x"C4DC0014";
end if;
if pc = 27664 then
	inst <= x"C49C000C";
end if;
if pc = 27668 then
	inst <= x"C17DFFFC";
end if;
if pc = 27672 then
	inst <= x"004A0000";
end if;
if pc = 27676 then
	inst <= x"002E0000";
end if;
if pc = 27680 then
	inst <= x"03DC0020";
end if;
if pc = 27684 then
	inst <= x"037E000C";
end if;
if pc = 27688 then
	inst <= x"C57DFFFC";
end if;
if pc = 27692 then
	inst <= x"82006424";
end if;
if pc = 27696 then
	inst <= x"07DC0020";
end if;
if pc = 27700 then
	inst <= x"C03C000C";
end if;
if pc = 27704 then
	inst <= x"C0420008";
end if;
if pc = 27708 then
	inst <= x"0260FFFF";
end if;
if pc = 27712 then
	inst <= x"82466CE8";
end if;
if pc = 27716 then
	inst <= x"22440220";
end if;
if pc = 27720 then
	inst <= x"C07C0014";
end if;
if pc = 27724 then
	inst <= x"D0464000";
end if;
if pc = 27728 then
	inst <= x"02800000";
end if;
if pc = 27732 then
	inst <= x"C0BC0000";
end if;
if pc = 27736 then
	inst <= x"C17DFFFC";
end if;
if pc = 27740 then
	inst <= x"006A0000";
end if;
if pc = 27744 then
	inst <= x"00280000";
end if;
if pc = 27748 then
	inst <= x"03DC0020";
end if;
if pc = 27752 then
	inst <= x"037E000C";
end if;
if pc = 27756 then
	inst <= x"C57DFFFC";
end if;
if pc = 27760 then
	inst <= x"82006424";
end if;
if pc = 27764 then
	inst <= x"07DC0020";
end if;
if pc = 27768 then
	inst <= x"C03C000C";
end if;
if pc = 27772 then
	inst <= x"C042000C";
end if;
if pc = 27776 then
	inst <= x"0260FFFF";
end if;
if pc = 27780 then
	inst <= x"82466CE4";
end if;
if pc = 27784 then
	inst <= x"22440220";
end if;
if pc = 27788 then
	inst <= x"C07C0014";
end if;
if pc = 27792 then
	inst <= x"D0464000";
end if;
if pc = 27796 then
	inst <= x"02600000";
end if;
if pc = 27800 then
	inst <= x"C09C0000";
end if;
if pc = 27804 then
	inst <= x"C17DFFFC";
end if;
if pc = 27808 then
	inst <= x"00260000";
end if;
if pc = 27812 then
	inst <= x"00680000";
end if;
if pc = 27816 then
	inst <= x"03DC0020";
end if;
if pc = 27820 then
	inst <= x"037E000C";
end if;
if pc = 27824 then
	inst <= x"C57DFFFC";
end if;
if pc = 27828 then
	inst <= x"82006424";
end if;
if pc = 27832 then
	inst <= x"07DC0020";
end if;
if pc = 27836 then
	inst <= x"02200004";
end if;
if pc = 27840 then
	inst <= x"C05C000C";
end if;
if pc = 27844 then
	inst <= x"C07C0000";
end if;
if pc = 27848 then
	inst <= x"C17DFFFC";
end if;
if pc = 27852 then
	inst <= x"03DC0020";
end if;
if pc = 27856 then
	inst <= x"037E000C";
end if;
if pc = 27860 then
	inst <= x"C57DFFFC";
end if;
if pc = 27864 then
	inst <= x"82006878";
end if;
if pc = 27868 then
	inst <= x"07DC0020";
end if;
if pc = 27872 then
	inst <= x"82006CE4";
end if;
if pc = 27876 then
	inst <= x"82006CE8";
end if;
if pc = 27880 then
	inst <= x"82006CEC";
end if;
if pc = 27884 then
	inst <= x"C03C0008";
end if;
if pc = 27888 then
	inst <= x"02220001";
end if;
if pc = 27892 then
	inst <= x"22420220";
end if;
if pc = 27896 then
	inst <= x"C07C0004";
end if;
if pc = 27900 then
	inst <= x"D0464000";
end if;
if pc = 27904 then
	inst <= x"C0840000";
end if;
if pc = 27908 then
	inst <= x"02A0FFFF";
end if;
if pc = 27912 then
	inst <= x"828A6F84";
end if;
if pc = 27916 then
	inst <= x"02A00063";
end if;
if pc = 27920 then
	inst <= x"C43C0018";
end if;
if pc = 27924 then
	inst <= x"828A6EB4";
end if;
if pc = 27928 then
	inst <= x"02A000C8";
end if;
if pc = 27932 then
	inst <= x"22C80220";
end if;
if pc = 27936 then
	inst <= x"D0AAC000";
end if;
if pc = 27940 then
	inst <= x"C0CA0028";
end if;
if pc = 27944 then
	inst <= x"C82C0000";
end if;
if pc = 27948 then
	inst <= x"C84C0004";
end if;
if pc = 27952 then
	inst <= x"C86C0008";
end if;
if pc = 27956 then
	inst <= x"C0FC0000";
end if;
if pc = 27960 then
	inst <= x"C10E0004";
end if;
if pc = 27964 then
	inst <= x"22880220";
end if;
if pc = 27968 then
	inst <= x"D0908000";
end if;
if pc = 27972 then
	inst <= x"C10A0004";
end if;
if pc = 27976 then
	inst <= x"03200001";
end if;
if pc = 27980 then
	inst <= x"C45C001C";
end if;
if pc = 27984 then
	inst <= x"83126DB0";
end if;
if pc = 27988 then
	inst <= x"03200002";
end if;
if pc = 27992 then
	inst <= x"83126D84";
end if;
if pc = 27996 then
	inst <= x"C17DFFFC";
end if;
if pc = 28000 then
	inst <= x"006C0000";
end if;
if pc = 28004 then
	inst <= x"00480000";
end if;
if pc = 28008 then
	inst <= x"002A0000";
end if;
if pc = 28012 then
	inst <= x"03DC0028";
end if;
if pc = 28016 then
	inst <= x"037E000C";
end if;
if pc = 28020 then
	inst <= x"C57DFFFC";
end if;
if pc = 28024 then
	inst <= x"82003BD4";
end if;
if pc = 28028 then
	inst <= x"07DC0028";
end if;
if pc = 28032 then
	inst <= x"82006DAC";
end if;
if pc = 28036 then
	inst <= x"C8280000";
end if;
if pc = 28040 then
	inst <= x"8E206D94";
end if;
if pc = 28044 then
	inst <= x"02200000";
end if;
if pc = 28048 then
	inst <= x"82006DAC";
end if;
if pc = 28052 then
	inst <= x"02A002AC";
end if;
if pc = 28056 then
	inst <= x"C8280000";
end if;
if pc = 28060 then
	inst <= x"C84C000C";
end if;
if pc = 28064 then
	inst <= x"48224000";
end if;
if pc = 28068 then
	inst <= x"CC2A0000";
end if;
if pc = 28072 then
	inst <= x"02200001";
end if;
if pc = 28076 then
	inst <= x"82006DD8";
end if;
if pc = 28080 then
	inst <= x"C0CE0000";
end if;
if pc = 28084 then
	inst <= x"C17DFFFC";
end if;
if pc = 28088 then
	inst <= x"00680000";
end if;
if pc = 28092 then
	inst <= x"004C0000";
end if;
if pc = 28096 then
	inst <= x"002A0000";
end if;
if pc = 28100 then
	inst <= x"03DC0028";
end if;
if pc = 28104 then
	inst <= x"037E000C";
end if;
if pc = 28108 then
	inst <= x"C57DFFFC";
end if;
if pc = 28112 then
	inst <= x"8200389C";
end if;
if pc = 28116 then
	inst <= x"07DC0028";
end if;
if pc = 28120 then
	inst <= x"82206EB0";
end if;
if pc = 28124 then
	inst <= x"022002AC";
end if;
if pc = 28128 then
	inst <= x"C8220000";
end if;
if pc = 28132 then
	inst <= x"022002B4";
end if;
if pc = 28136 then
	inst <= x"C8420000";
end if;
if pc = 28140 then
	inst <= x"8E246DF4";
end if;
if pc = 28144 then
	inst <= x"82006EAC";
end if;
if pc = 28148 then
	inst <= x"C03C001C";
end if;
if pc = 28152 then
	inst <= x"C0420004";
end if;
if pc = 28156 then
	inst <= x"0260FFFF";
end if;
if pc = 28160 then
	inst <= x"82466EAC";
end if;
if pc = 28164 then
	inst <= x"026001E0";
end if;
if pc = 28168 then
	inst <= x"22440220";
end if;
if pc = 28172 then
	inst <= x"D0464000";
end if;
if pc = 28176 then
	inst <= x"02800000";
end if;
if pc = 28180 then
	inst <= x"C0BC0000";
end if;
if pc = 28184 then
	inst <= x"C47C0020";
end if;
if pc = 28188 then
	inst <= x"C17DFFFC";
end if;
if pc = 28192 then
	inst <= x"006A0000";
end if;
if pc = 28196 then
	inst <= x"00280000";
end if;
if pc = 28200 then
	inst <= x"03DC002C";
end if;
if pc = 28204 then
	inst <= x"037E000C";
end if;
if pc = 28208 then
	inst <= x"C57DFFFC";
end if;
if pc = 28212 then
	inst <= x"82006424";
end if;
if pc = 28216 then
	inst <= x"07DC002C";
end if;
if pc = 28220 then
	inst <= x"C03C001C";
end if;
if pc = 28224 then
	inst <= x"C0420008";
end if;
if pc = 28228 then
	inst <= x"0260FFFF";
end if;
if pc = 28232 then
	inst <= x"82466EA8";
end if;
if pc = 28236 then
	inst <= x"22440220";
end if;
if pc = 28240 then
	inst <= x"C07C0020";
end if;
if pc = 28244 then
	inst <= x"D0464000";
end if;
if pc = 28248 then
	inst <= x"02600000";
end if;
if pc = 28252 then
	inst <= x"C09C0000";
end if;
if pc = 28256 then
	inst <= x"C17DFFFC";
end if;
if pc = 28260 then
	inst <= x"00260000";
end if;
if pc = 28264 then
	inst <= x"00680000";
end if;
if pc = 28268 then
	inst <= x"03DC002C";
end if;
if pc = 28272 then
	inst <= x"037E000C";
end if;
if pc = 28276 then
	inst <= x"C57DFFFC";
end if;
if pc = 28280 then
	inst <= x"82006424";
end if;
if pc = 28284 then
	inst <= x"07DC002C";
end if;
if pc = 28288 then
	inst <= x"02200003";
end if;
if pc = 28292 then
	inst <= x"C05C001C";
end if;
if pc = 28296 then
	inst <= x"C07C0000";
end if;
if pc = 28300 then
	inst <= x"C17DFFFC";
end if;
if pc = 28304 then
	inst <= x"03DC002C";
end if;
if pc = 28308 then
	inst <= x"037E000C";
end if;
if pc = 28312 then
	inst <= x"C57DFFFC";
end if;
if pc = 28316 then
	inst <= x"82006878";
end if;
if pc = 28320 then
	inst <= x"07DC002C";
end if;
if pc = 28324 then
	inst <= x"82006EA8";
end if;
if pc = 28328 then
	inst <= x"82006EAC";
end if;
if pc = 28332 then
	inst <= x"82006EB0";
end if;
if pc = 28336 then
	inst <= x"82006F70";
end if;
if pc = 28340 then
	inst <= x"C0840004";
end if;
if pc = 28344 then
	inst <= x"02A0FFFF";
end if;
if pc = 28348 then
	inst <= x"828A6F70";
end if;
if pc = 28352 then
	inst <= x"02A001E0";
end if;
if pc = 28356 then
	inst <= x"22880220";
end if;
if pc = 28360 then
	inst <= x"D08A8000";
end if;
if pc = 28364 then
	inst <= x"02C00000";
end if;
if pc = 28368 then
	inst <= x"C0FC0000";
end if;
if pc = 28372 then
	inst <= x"C4BC0024";
end if;
if pc = 28376 then
	inst <= x"C45C001C";
end if;
if pc = 28380 then
	inst <= x"C17DFFFC";
end if;
if pc = 28384 then
	inst <= x"006E0000";
end if;
if pc = 28388 then
	inst <= x"00480000";
end if;
if pc = 28392 then
	inst <= x"002C0000";
end if;
if pc = 28396 then
	inst <= x"03DC0030";
end if;
if pc = 28400 then
	inst <= x"037E000C";
end if;
if pc = 28404 then
	inst <= x"C57DFFFC";
end if;
if pc = 28408 then
	inst <= x"82006424";
end if;
if pc = 28412 then
	inst <= x"07DC0030";
end if;
if pc = 28416 then
	inst <= x"C03C001C";
end if;
if pc = 28420 then
	inst <= x"C0420008";
end if;
if pc = 28424 then
	inst <= x"0260FFFF";
end if;
if pc = 28428 then
	inst <= x"82466F6C";
end if;
if pc = 28432 then
	inst <= x"22440220";
end if;
if pc = 28436 then
	inst <= x"C07C0024";
end if;
if pc = 28440 then
	inst <= x"D0464000";
end if;
if pc = 28444 then
	inst <= x"02600000";
end if;
if pc = 28448 then
	inst <= x"C09C0000";
end if;
if pc = 28452 then
	inst <= x"C17DFFFC";
end if;
if pc = 28456 then
	inst <= x"00260000";
end if;
if pc = 28460 then
	inst <= x"00680000";
end if;
if pc = 28464 then
	inst <= x"03DC0030";
end if;
if pc = 28468 then
	inst <= x"037E000C";
end if;
if pc = 28472 then
	inst <= x"C57DFFFC";
end if;
if pc = 28476 then
	inst <= x"82006424";
end if;
if pc = 28480 then
	inst <= x"07DC0030";
end if;
if pc = 28484 then
	inst <= x"02200003";
end if;
if pc = 28488 then
	inst <= x"C05C001C";
end if;
if pc = 28492 then
	inst <= x"C07C0000";
end if;
if pc = 28496 then
	inst <= x"C17DFFFC";
end if;
if pc = 28500 then
	inst <= x"03DC0030";
end if;
if pc = 28504 then
	inst <= x"037E000C";
end if;
if pc = 28508 then
	inst <= x"C57DFFFC";
end if;
if pc = 28512 then
	inst <= x"82006878";
end if;
if pc = 28516 then
	inst <= x"07DC0030";
end if;
if pc = 28520 then
	inst <= x"82006F6C";
end if;
if pc = 28524 then
	inst <= x"82006F70";
end if;
if pc = 28528 then
	inst <= x"C03C0018";
end if;
if pc = 28532 then
	inst <= x"02220001";
end if;
if pc = 28536 then
	inst <= x"C05C0004";
end if;
if pc = 28540 then
	inst <= x"C07C0000";
end if;
if pc = 28544 then
	inst <= x"820069E8";
end if;
if pc = 28548 then
	inst <= x"C1FDFFFC";
end if;
if pc = 28552 then
	inst <= x"C1FDFFFC";
end if;
if pc = 28556 then
	inst <= x"024002B8";
end if;
if pc = 28560 then
	inst <= x"C8240000";
end if;
if pc = 28564 then
	inst <= x"C0620014";
end if;
if pc = 28568 then
	inst <= x"C8460000";
end if;
if pc = 28572 then
	inst <= x"44224000";
end if;
if pc = 28576 then
	inst <= x"C8440004";
end if;
if pc = 28580 then
	inst <= x"C0620014";
end if;
if pc = 28584 then
	inst <= x"C8660004";
end if;
if pc = 28588 then
	inst <= x"44446000";
end if;
if pc = 28592 then
	inst <= x"C8640008";
end if;
if pc = 28596 then
	inst <= x"C0420014";
end if;
if pc = 28600 then
	inst <= x"C8840008";
end if;
if pc = 28604 then
	inst <= x"44668000";
end if;
if pc = 28608 then
	inst <= x"C0420010";
end if;
if pc = 28612 then
	inst <= x"C8840000";
end if;
if pc = 28616 then
	inst <= x"48828000";
end if;
if pc = 28620 then
	inst <= x"C0420010";
end if;
if pc = 28624 then
	inst <= x"C8A40004";
end if;
if pc = 28628 then
	inst <= x"48A4A000";
end if;
if pc = 28632 then
	inst <= x"C0420010";
end if;
if pc = 28636 then
	inst <= x"C8C40008";
end if;
if pc = 28640 then
	inst <= x"48C6C000";
end if;
if pc = 28644 then
	inst <= x"C042000C";
end if;
if pc = 28648 then
	inst <= x"C43C0000";
end if;
if pc = 28652 then
	inst <= x"82407138";
end if;
if pc = 28656 then
	inst <= x"024002C8";
end if;
if pc = 28660 then
	inst <= x"C0620024";
end if;
if pc = 28664 then
	inst <= x"C8E60008";
end if;
if pc = 28668 then
	inst <= x"48E4E000";
end if;
if pc = 28672 then
	inst <= x"C0620024";
end if;
if pc = 28676 then
	inst <= x"C9060004";
end if;
if pc = 28680 then
	inst <= x"49070000";
end if;
if pc = 28684 then
	inst <= x"40EF0000";
end if;
if pc = 28688 then
	inst <= x"C9000080";
end if;
if pc = 28692 then
	inst <= x"CCDC0008";
end if;
if pc = 28696 then
	inst <= x"CC5C0010";
end if;
if pc = 28700 then
	inst <= x"CCBC0018";
end if;
if pc = 28704 then
	inst <= x"CD1C0020";
end if;
if pc = 28708 then
	inst <= x"CC7C0028";
end if;
if pc = 28712 then
	inst <= x"CC3C0030";
end if;
if pc = 28716 then
	inst <= x"C45C0038";
end if;
if pc = 28720 then
	inst <= x"CC9C0040";
end if;
if pc = 28724 then
	inst <= x"CCFC0048";
end if;
if pc = 28728 then
	inst <= x"C17DFFFC";
end if;
if pc = 28732 then
	inst <= x"40210000";
end if;
if pc = 28736 then
	inst <= x"03DC0058";
end if;
if pc = 28740 then
	inst <= x"037E000C";
end if;
if pc = 28744 then
	inst <= x"C57DFFFC";
end if;
if pc = 28748 then
	inst <= x"82000844";
end if;
if pc = 28752 then
	inst <= x"07DC0058";
end if;
if pc = 28756 then
	inst <= x"C85C0048";
end if;
if pc = 28760 then
	inst <= x"48242000";
end if;
if pc = 28764 then
	inst <= x"C85C0040";
end if;
if pc = 28768 then
	inst <= x"40242000";
end if;
if pc = 28772 then
	inst <= x"C03C0038";
end if;
if pc = 28776 then
	inst <= x"CC220000";
end if;
if pc = 28780 then
	inst <= x"C05C0000";
end if;
if pc = 28784 then
	inst <= x"C0640024";
end if;
if pc = 28788 then
	inst <= x"C8260008";
end if;
if pc = 28792 then
	inst <= x"C85C0030";
end if;
if pc = 28796 then
	inst <= x"48242000";
end if;
if pc = 28800 then
	inst <= x"C0640024";
end if;
if pc = 28804 then
	inst <= x"C8660000";
end if;
if pc = 28808 then
	inst <= x"C89C0028";
end if;
if pc = 28812 then
	inst <= x"48686000";
end if;
if pc = 28816 then
	inst <= x"40226000";
end if;
if pc = 28820 then
	inst <= x"C87C0020";
end if;
if pc = 28824 then
	inst <= x"CC3C0050";
end if;
if pc = 28828 then
	inst <= x"C17DFFFC";
end if;
if pc = 28832 then
	inst <= x"40206000";
end if;
if pc = 28836 then
	inst <= x"03DC0060";
end if;
if pc = 28840 then
	inst <= x"037E000C";
end if;
if pc = 28844 then
	inst <= x"C57DFFFC";
end if;
if pc = 28848 then
	inst <= x"82000844";
end if;
if pc = 28852 then
	inst <= x"07DC0060";
end if;
if pc = 28856 then
	inst <= x"C85C0050";
end if;
if pc = 28860 then
	inst <= x"48242000";
end if;
if pc = 28864 then
	inst <= x"C85C0018";
end if;
if pc = 28868 then
	inst <= x"40242000";
end if;
if pc = 28872 then
	inst <= x"C03C0038";
end if;
if pc = 28876 then
	inst <= x"CC220004";
end if;
if pc = 28880 then
	inst <= x"C05C0000";
end if;
if pc = 28884 then
	inst <= x"C0640024";
end if;
if pc = 28888 then
	inst <= x"C8260004";
end if;
if pc = 28892 then
	inst <= x"C85C0030";
end if;
if pc = 28896 then
	inst <= x"48242000";
end if;
if pc = 28900 then
	inst <= x"C0640024";
end if;
if pc = 28904 then
	inst <= x"C8460000";
end if;
if pc = 28908 then
	inst <= x"C87C0010";
end if;
if pc = 28912 then
	inst <= x"48464000";
end if;
if pc = 28916 then
	inst <= x"40224000";
end if;
if pc = 28920 then
	inst <= x"C85C0020";
end if;
if pc = 28924 then
	inst <= x"CC3C0058";
end if;
if pc = 28928 then
	inst <= x"C17DFFFC";
end if;
if pc = 28932 then
	inst <= x"40204000";
end if;
if pc = 28936 then
	inst <= x"03DC0068";
end if;
if pc = 28940 then
	inst <= x"037E000C";
end if;
if pc = 28944 then
	inst <= x"C57DFFFC";
end if;
if pc = 28948 then
	inst <= x"82000844";
end if;
if pc = 28952 then
	inst <= x"07DC0068";
end if;
if pc = 28956 then
	inst <= x"C85C0058";
end if;
if pc = 28960 then
	inst <= x"48242000";
end if;
if pc = 28964 then
	inst <= x"C85C0008";
end if;
if pc = 28968 then
	inst <= x"40242000";
end if;
if pc = 28972 then
	inst <= x"C03C0038";
end if;
if pc = 28976 then
	inst <= x"CC220008";
end if;
if pc = 28980 then
	inst <= x"82007148";
end if;
if pc = 28984 then
	inst <= x"024002C8";
end if;
if pc = 28988 then
	inst <= x"CC840000";
end if;
if pc = 28992 then
	inst <= x"CCA40004";
end if;
if pc = 28996 then
	inst <= x"CCC40008";
end if;
if pc = 29000 then
	inst <= x"022002C8";
end if;
if pc = 29004 then
	inst <= x"C05C0000";
end if;
if pc = 29008 then
	inst <= x"C0440018";
end if;
if pc = 29012 then
	inst <= x"8200161C";
end if;
if pc = 29016 then
	inst <= x"C0620000";
end if;
if pc = 29020 then
	inst <= x"028002D4";
end if;
if pc = 29024 then
	inst <= x"C0A20020";
end if;
if pc = 29028 then
	inst <= x"C82A0000";
end if;
if pc = 29032 then
	inst <= x"CC280000";
end if;
if pc = 29036 then
	inst <= x"C0A20020";
end if;
if pc = 29040 then
	inst <= x"C82A0004";
end if;
if pc = 29044 then
	inst <= x"CC280004";
end if;
if pc = 29048 then
	inst <= x"C0A20020";
end if;
if pc = 29052 then
	inst <= x"C82A0008";
end if;
if pc = 29056 then
	inst <= x"CC280008";
end if;
if pc = 29060 then
	inst <= x"02A00001";
end if;
if pc = 29064 then
	inst <= x"826A7710";
end if;
if pc = 29068 then
	inst <= x"02A00002";
end if;
if pc = 29072 then
	inst <= x"826A7648";
end if;
if pc = 29076 then
	inst <= x"02A00003";
end if;
if pc = 29080 then
	inst <= x"826A74E8";
end if;
if pc = 29084 then
	inst <= x"02A00004";
end if;
if pc = 29088 then
	inst <= x"826A71A8";
end if;
if pc = 29092 then
	inst <= x"C1FDFFFC";
end if;
if pc = 29096 then
	inst <= x"C8240000";
end if;
if pc = 29100 then
	inst <= x"C0620014";
end if;
if pc = 29104 then
	inst <= x"C8460000";
end if;
if pc = 29108 then
	inst <= x"44224000";
end if;
if pc = 29112 then
	inst <= x"C0620010";
end if;
if pc = 29116 then
	inst <= x"C8460000";
end if;
if pc = 29120 then
	inst <= x"C49C0000";
end if;
if pc = 29124 then
	inst <= x"C43C0004";
end if;
if pc = 29128 then
	inst <= x"C45C0008";
end if;
if pc = 29132 then
	inst <= x"CC3C0010";
end if;
if pc = 29136 then
	inst <= x"C17DFFFC";
end if;
if pc = 29140 then
	inst <= x"40204000";
end if;
if pc = 29144 then
	inst <= x"03DC0020";
end if;
if pc = 29148 then
	inst <= x"037E000C";
end if;
if pc = 29152 then
	inst <= x"C57DFFFC";
end if;
if pc = 29156 then
	inst <= x"8200083C";
end if;
if pc = 29160 then
	inst <= x"07DC0020";
end if;
if pc = 29164 then
	inst <= x"C85C0010";
end if;
if pc = 29168 then
	inst <= x"48242000";
end if;
if pc = 29172 then
	inst <= x"C03C0008";
end if;
if pc = 29176 then
	inst <= x"C8420008";
end if;
if pc = 29180 then
	inst <= x"C05C0004";
end if;
if pc = 29184 then
	inst <= x"C0640014";
end if;
if pc = 29188 then
	inst <= x"C8660008";
end if;
if pc = 29192 then
	inst <= x"44446000";
end if;
if pc = 29196 then
	inst <= x"C0640010";
end if;
if pc = 29200 then
	inst <= x"C8660008";
end if;
if pc = 29204 then
	inst <= x"CC3C0018";
end if;
if pc = 29208 then
	inst <= x"CC5C0020";
end if;
if pc = 29212 then
	inst <= x"C17DFFFC";
end if;
if pc = 29216 then
	inst <= x"40206000";
end if;
if pc = 29220 then
	inst <= x"03DC0030";
end if;
if pc = 29224 then
	inst <= x"037E000C";
end if;
if pc = 29228 then
	inst <= x"C57DFFFC";
end if;
if pc = 29232 then
	inst <= x"8200083C";
end if;
if pc = 29236 then
	inst <= x"07DC0030";
end if;
if pc = 29240 then
	inst <= x"C85C0020";
end if;
if pc = 29244 then
	inst <= x"48242000";
end if;
if pc = 29248 then
	inst <= x"C85C0018";
end if;
if pc = 29252 then
	inst <= x"48644000";
end if;
if pc = 29256 then
	inst <= x"48822000";
end if;
if pc = 29260 then
	inst <= x"40668000";
end if;
if pc = 29264 then
	inst <= x"8E40725C";
end if;
if pc = 29268 then
	inst <= x"40804000";
end if;
if pc = 29272 then
	inst <= x"82007260";
end if;
if pc = 29276 then
	inst <= x"44804000";
end if;
if pc = 29280 then
	inst <= x"C8A0006C";
end if;
if pc = 29284 then
	inst <= x"CCBC0028";
end if;
if pc = 29288 then
	inst <= x"CC7C0030";
end if;
if pc = 29292 then
	inst <= x"8E8A7310";
end if;
if pc = 29296 then
	inst <= x"CC3C0038";
end if;
if pc = 29300 then
	inst <= x"C17DFFFC";
end if;
if pc = 29304 then
	inst <= x"40204000";
end if;
if pc = 29308 then
	inst <= x"03DC0048";
end if;
if pc = 29312 then
	inst <= x"037E000C";
end if;
if pc = 29316 then
	inst <= x"C57DFFFC";
end if;
if pc = 29320 then
	inst <= x"82000844";
end if;
if pc = 29324 then
	inst <= x"07DC0048";
end if;
if pc = 29328 then
	inst <= x"C85C0038";
end if;
if pc = 29332 then
	inst <= x"48242000";
end if;
if pc = 29336 then
	inst <= x"8E2072A0";
end if;
if pc = 29340 then
	inst <= x"820072A4";
end if;
if pc = 29344 then
	inst <= x"44202000";
end if;
if pc = 29348 then
	inst <= x"C8400068";
end if;
if pc = 29352 then
	inst <= x"48442000";
end if;
if pc = 29356 then
	inst <= x"C8600064";
end if;
if pc = 29360 then
	inst <= x"44446000";
end if;
if pc = 29364 then
	inst <= x"48442000";
end if;
if pc = 29368 then
	inst <= x"C8600060";
end if;
if pc = 29372 then
	inst <= x"44446000";
end if;
if pc = 29376 then
	inst <= x"48442000";
end if;
if pc = 29380 then
	inst <= x"C860005C";
end if;
if pc = 29384 then
	inst <= x"40446000";
end if;
if pc = 29388 then
	inst <= x"48242000";
end if;
if pc = 29392 then
	inst <= x"C8400058";
end if;
if pc = 29396 then
	inst <= x"44224000";
end if;
if pc = 29400 then
	inst <= x"C8400054";
end if;
if pc = 29404 then
	inst <= x"48224000";
end if;
if pc = 29408 then
	inst <= x"C8400050";
end if;
if pc = 29412 then
	inst <= x"CC3C0040";
end if;
if pc = 29416 then
	inst <= x"C17DFFFC";
end if;
if pc = 29420 then
	inst <= x"40204000";
end if;
if pc = 29424 then
	inst <= x"03DC0050";
end if;
if pc = 29428 then
	inst <= x"037E000C";
end if;
if pc = 29432 then
	inst <= x"C57DFFFC";
end if;
if pc = 29436 then
	inst <= x"82000844";
end if;
if pc = 29440 then
	inst <= x"07DC0050";
end if;
if pc = 29444 then
	inst <= x"C85C0040";
end if;
if pc = 29448 then
	inst <= x"48242000";
end if;
if pc = 29452 then
	inst <= x"82007314";
end if;
if pc = 29456 then
	inst <= x"C820004C";
end if;
if pc = 29460 then
	inst <= x"54220000";
end if;
if pc = 29464 then
	inst <= x"8E027338";
end if;
if pc = 29468 then
	inst <= x"58420000";
end if;
if pc = 29472 then
	inst <= x"8A427330";
end if;
if pc = 29476 then
	inst <= x"06220001";
end if;
if pc = 29480 then
	inst <= x"58420000";
end if;
if pc = 29484 then
	inst <= x"82007334";
end if;
if pc = 29488 then
	inst <= x"40402000";
end if;
if pc = 29492 then
	inst <= x"8200733C";
end if;
if pc = 29496 then
	inst <= x"58420000";
end if;
if pc = 29500 then
	inst <= x"44224000";
end if;
if pc = 29504 then
	inst <= x"C03C0008";
end if;
if pc = 29508 then
	inst <= x"C8420004";
end if;
if pc = 29512 then
	inst <= x"C03C0004";
end if;
if pc = 29516 then
	inst <= x"C0420014";
end if;
if pc = 29520 then
	inst <= x"C8640004";
end if;
if pc = 29524 then
	inst <= x"44446000";
end if;
if pc = 29528 then
	inst <= x"C0220010";
end if;
if pc = 29532 then
	inst <= x"C8620004";
end if;
if pc = 29536 then
	inst <= x"CC3C0048";
end if;
if pc = 29540 then
	inst <= x"CC5C0050";
end if;
if pc = 29544 then
	inst <= x"C17DFFFC";
end if;
if pc = 29548 then
	inst <= x"40206000";
end if;
if pc = 29552 then
	inst <= x"03DC0060";
end if;
if pc = 29556 then
	inst <= x"037E000C";
end if;
if pc = 29560 then
	inst <= x"C57DFFFC";
end if;
if pc = 29564 then
	inst <= x"8200083C";
end if;
if pc = 29568 then
	inst <= x"07DC0060";
end if;
if pc = 29572 then
	inst <= x"C85C0050";
end if;
if pc = 29576 then
	inst <= x"48242000";
end if;
if pc = 29580 then
	inst <= x"C85C0030";
end if;
if pc = 29584 then
	inst <= x"8E40739C";
end if;
if pc = 29588 then
	inst <= x"40604000";
end if;
if pc = 29592 then
	inst <= x"820073A0";
end if;
if pc = 29596 then
	inst <= x"44604000";
end if;
if pc = 29600 then
	inst <= x"C89C0028";
end if;
if pc = 29604 then
	inst <= x"8E687448";
end if;
if pc = 29608 then
	inst <= x"CC3C0058";
end if;
if pc = 29612 then
	inst <= x"C17DFFFC";
end if;
if pc = 29616 then
	inst <= x"40204000";
end if;
if pc = 29620 then
	inst <= x"03DC0068";
end if;
if pc = 29624 then
	inst <= x"037E000C";
end if;
if pc = 29628 then
	inst <= x"C57DFFFC";
end if;
if pc = 29632 then
	inst <= x"82000844";
end if;
if pc = 29636 then
	inst <= x"07DC0068";
end if;
if pc = 29640 then
	inst <= x"C85C0058";
end if;
if pc = 29644 then
	inst <= x"48242000";
end if;
if pc = 29648 then
	inst <= x"8E2073D8";
end if;
if pc = 29652 then
	inst <= x"820073DC";
end if;
if pc = 29656 then
	inst <= x"44202000";
end if;
if pc = 29660 then
	inst <= x"C8400068";
end if;
if pc = 29664 then
	inst <= x"48442000";
end if;
if pc = 29668 then
	inst <= x"C8600064";
end if;
if pc = 29672 then
	inst <= x"44446000";
end if;
if pc = 29676 then
	inst <= x"48442000";
end if;
if pc = 29680 then
	inst <= x"C8600060";
end if;
if pc = 29684 then
	inst <= x"44446000";
end if;
if pc = 29688 then
	inst <= x"48442000";
end if;
if pc = 29692 then
	inst <= x"C860005C";
end if;
if pc = 29696 then
	inst <= x"40446000";
end if;
if pc = 29700 then
	inst <= x"48242000";
end if;
if pc = 29704 then
	inst <= x"C8400058";
end if;
if pc = 29708 then
	inst <= x"44224000";
end if;
if pc = 29712 then
	inst <= x"C8400054";
end if;
if pc = 29716 then
	inst <= x"48224000";
end if;
if pc = 29720 then
	inst <= x"C8400050";
end if;
if pc = 29724 then
	inst <= x"CC3C0060";
end if;
if pc = 29728 then
	inst <= x"C17DFFFC";
end if;
if pc = 29732 then
	inst <= x"40204000";
end if;
if pc = 29736 then
	inst <= x"03DC0070";
end if;
if pc = 29740 then
	inst <= x"037E000C";
end if;
if pc = 29744 then
	inst <= x"C57DFFFC";
end if;
if pc = 29748 then
	inst <= x"82000844";
end if;
if pc = 29752 then
	inst <= x"07DC0070";
end if;
if pc = 29756 then
	inst <= x"C85C0060";
end if;
if pc = 29760 then
	inst <= x"48242000";
end if;
if pc = 29764 then
	inst <= x"8200744C";
end if;
if pc = 29768 then
	inst <= x"C820004C";
end if;
if pc = 29772 then
	inst <= x"54220000";
end if;
if pc = 29776 then
	inst <= x"8E027470";
end if;
if pc = 29780 then
	inst <= x"58420000";
end if;
if pc = 29784 then
	inst <= x"8A427468";
end if;
if pc = 29788 then
	inst <= x"06220001";
end if;
if pc = 29792 then
	inst <= x"58420000";
end if;
if pc = 29796 then
	inst <= x"8200746C";
end if;
if pc = 29800 then
	inst <= x"40402000";
end if;
if pc = 29804 then
	inst <= x"82007474";
end if;
if pc = 29808 then
	inst <= x"58420000";
end if;
if pc = 29812 then
	inst <= x"44224000";
end if;
if pc = 29816 then
	inst <= x"C8400048";
end if;
if pc = 29820 then
	inst <= x"C86000A4";
end if;
if pc = 29824 then
	inst <= x"C89C0048";
end if;
if pc = 29828 then
	inst <= x"44868000";
end if;
if pc = 29832 then
	inst <= x"48888000";
end if;
if pc = 29836 then
	inst <= x"44448000";
end if;
if pc = 29840 then
	inst <= x"44262000";
end if;
if pc = 29844 then
	inst <= x"48222000";
end if;
if pc = 29848 then
	inst <= x"44242000";
end if;
if pc = 29852 then
	inst <= x"8E2074A4";
end if;
if pc = 29856 then
	inst <= x"820074A8";
end if;
if pc = 29860 then
	inst <= x"40200000";
end if;
if pc = 29864 then
	inst <= x"C8400044";
end if;
if pc = 29868 then
	inst <= x"48242000";
end if;
if pc = 29872 then
	inst <= x"C8400040";
end if;
if pc = 29876 then
	inst <= x"CC3C0068";
end if;
if pc = 29880 then
	inst <= x"C17DFFFC";
end if;
if pc = 29884 then
	inst <= x"40204000";
end if;
if pc = 29888 then
	inst <= x"03DC0078";
end if;
if pc = 29892 then
	inst <= x"037E000C";
end if;
if pc = 29896 then
	inst <= x"C57DFFFC";
end if;
if pc = 29900 then
	inst <= x"82000844";
end if;
if pc = 29904 then
	inst <= x"07DC0078";
end if;
if pc = 29908 then
	inst <= x"C85C0068";
end if;
if pc = 29912 then
	inst <= x"48242000";
end if;
if pc = 29916 then
	inst <= x"C03C0000";
end if;
if pc = 29920 then
	inst <= x"CC220008";
end if;
if pc = 29924 then
	inst <= x"C1FDFFFC";
end if;
if pc = 29928 then
	inst <= x"C8240000";
end if;
if pc = 29932 then
	inst <= x"C0620014";
end if;
if pc = 29936 then
	inst <= x"C8460000";
end if;
if pc = 29940 then
	inst <= x"44224000";
end if;
if pc = 29944 then
	inst <= x"C8440008";
end if;
if pc = 29948 then
	inst <= x"C0220014";
end if;
if pc = 29952 then
	inst <= x"C8620008";
end if;
if pc = 29956 then
	inst <= x"44446000";
end if;
if pc = 29960 then
	inst <= x"48222000";
end if;
if pc = 29964 then
	inst <= x"48444000";
end if;
if pc = 29968 then
	inst <= x"40224000";
end if;
if pc = 29972 then
	inst <= x"C49C0000";
end if;
if pc = 29976 then
	inst <= x"C17DFFFC";
end if;
if pc = 29980 then
	inst <= x"03DC0078";
end if;
if pc = 29984 then
	inst <= x"037E000C";
end if;
if pc = 29988 then
	inst <= x"C57DFFFC";
end if;
if pc = 29992 then
	inst <= x"8200083C";
end if;
if pc = 29996 then
	inst <= x"07DC0078";
end if;
if pc = 30000 then
	inst <= x"C840003C";
end if;
if pc = 30004 then
	inst <= x"CC3C0070";
end if;
if pc = 30008 then
	inst <= x"C17DFFFC";
end if;
if pc = 30012 then
	inst <= x"40204000";
end if;
if pc = 30016 then
	inst <= x"03DC0080";
end if;
if pc = 30020 then
	inst <= x"037E000C";
end if;
if pc = 30024 then
	inst <= x"C57DFFFC";
end if;
if pc = 30028 then
	inst <= x"82000844";
end if;
if pc = 30032 then
	inst <= x"07DC0080";
end if;
if pc = 30036 then
	inst <= x"C85C0070";
end if;
if pc = 30040 then
	inst <= x"48242000";
end if;
if pc = 30044 then
	inst <= x"54220000";
end if;
if pc = 30048 then
	inst <= x"8E027580";
end if;
if pc = 30052 then
	inst <= x"58420000";
end if;
if pc = 30056 then
	inst <= x"8A427578";
end if;
if pc = 30060 then
	inst <= x"06220001";
end if;
if pc = 30064 then
	inst <= x"58420000";
end if;
if pc = 30068 then
	inst <= x"8200757C";
end if;
if pc = 30072 then
	inst <= x"40402000";
end if;
if pc = 30076 then
	inst <= x"82007584";
end if;
if pc = 30080 then
	inst <= x"58420000";
end if;
if pc = 30084 then
	inst <= x"44224000";
end if;
if pc = 30088 then
	inst <= x"C8400050";
end if;
if pc = 30092 then
	inst <= x"48224000";
end if;
if pc = 30096 then
	inst <= x"C8400098";
end if;
if pc = 30100 then
	inst <= x"8E2475B8";
end if;
if pc = 30104 then
	inst <= x"44224000";
end if;
if pc = 30108 then
	inst <= x"C17DFFFC";
end if;
if pc = 30112 then
	inst <= x"03DC0080";
end if;
if pc = 30116 then
	inst <= x"037E000C";
end if;
if pc = 30120 then
	inst <= x"C57DFFFC";
end if;
if pc = 30124 then
	inst <= x"82001270";
end if;
if pc = 30128 then
	inst <= x"07DC0080";
end if;
if pc = 30132 then
	inst <= x"82007620";
end if;
if pc = 30136 then
	inst <= x"8E027604";
end if;
if pc = 30140 then
	inst <= x"C8600090";
end if;
if pc = 30144 then
	inst <= x"8E6275E4";
end if;
if pc = 30148 then
	inst <= x"40224000";
end if;
if pc = 30152 then
	inst <= x"C17DFFFC";
end if;
if pc = 30156 then
	inst <= x"03DC0080";
end if;
if pc = 30160 then
	inst <= x"037E000C";
end if;
if pc = 30164 then
	inst <= x"C57DFFFC";
end if;
if pc = 30168 then
	inst <= x"82001270";
end if;
if pc = 30172 then
	inst <= x"07DC0080";
end if;
if pc = 30176 then
	inst <= x"82007600";
end if;
if pc = 30180 then
	inst <= x"02200001";
end if;
if pc = 30184 then
	inst <= x"C17DFFFC";
end if;
if pc = 30188 then
	inst <= x"03DC0080";
end if;
if pc = 30192 then
	inst <= x"037E000C";
end if;
if pc = 30196 then
	inst <= x"C57DFFFC";
end if;
if pc = 30200 then
	inst <= x"82000B88";
end if;
if pc = 30204 then
	inst <= x"07DC0080";
end if;
if pc = 30208 then
	inst <= x"82007620";
end if;
if pc = 30212 then
	inst <= x"0220FFFF";
end if;
if pc = 30216 then
	inst <= x"C17DFFFC";
end if;
if pc = 30220 then
	inst <= x"03DC0080";
end if;
if pc = 30224 then
	inst <= x"037E000C";
end if;
if pc = 30228 then
	inst <= x"C57DFFFC";
end if;
if pc = 30232 then
	inst <= x"82000B88";
end if;
if pc = 30236 then
	inst <= x"07DC0080";
end if;
if pc = 30240 then
	inst <= x"48222000";
end if;
if pc = 30244 then
	inst <= x"C8400044";
end if;
if pc = 30248 then
	inst <= x"48624000";
end if;
if pc = 30252 then
	inst <= x"C03C0000";
end if;
if pc = 30256 then
	inst <= x"CC620004";
end if;
if pc = 30260 then
	inst <= x"C86000A8";
end if;
if pc = 30264 then
	inst <= x"44262000";
end if;
if pc = 30268 then
	inst <= x"48224000";
end if;
if pc = 30272 then
	inst <= x"CC220008";
end if;
if pc = 30276 then
	inst <= x"C1FDFFFC";
end if;
if pc = 30280 then
	inst <= x"C8240004";
end if;
if pc = 30284 then
	inst <= x"C8400038";
end if;
if pc = 30288 then
	inst <= x"48224000";
end if;
if pc = 30292 then
	inst <= x"C8400098";
end if;
if pc = 30296 then
	inst <= x"C49C0000";
end if;
if pc = 30300 then
	inst <= x"8E247680";
end if;
if pc = 30304 then
	inst <= x"44224000";
end if;
if pc = 30308 then
	inst <= x"C17DFFFC";
end if;
if pc = 30312 then
	inst <= x"03DC0080";
end if;
if pc = 30316 then
	inst <= x"037E000C";
end if;
if pc = 30320 then
	inst <= x"C57DFFFC";
end if;
if pc = 30324 then
	inst <= x"82000EC4";
end if;
if pc = 30328 then
	inst <= x"07DC0080";
end if;
if pc = 30332 then
	inst <= x"820076E8";
end if;
if pc = 30336 then
	inst <= x"8E0276CC";
end if;
if pc = 30340 then
	inst <= x"C8600090";
end if;
if pc = 30344 then
	inst <= x"8E6276AC";
end if;
if pc = 30348 then
	inst <= x"40224000";
end if;
if pc = 30352 then
	inst <= x"C17DFFFC";
end if;
if pc = 30356 then
	inst <= x"03DC0080";
end if;
if pc = 30360 then
	inst <= x"037E000C";
end if;
if pc = 30364 then
	inst <= x"C57DFFFC";
end if;
if pc = 30368 then
	inst <= x"82000EC4";
end if;
if pc = 30372 then
	inst <= x"07DC0080";
end if;
if pc = 30376 then
	inst <= x"820076C8";
end if;
if pc = 30380 then
	inst <= x"02200001";
end if;
if pc = 30384 then
	inst <= x"C17DFFFC";
end if;
if pc = 30388 then
	inst <= x"03DC0080";
end if;
if pc = 30392 then
	inst <= x"037E000C";
end if;
if pc = 30396 then
	inst <= x"C57DFFFC";
end if;
if pc = 30400 then
	inst <= x"8200084C";
end if;
if pc = 30404 then
	inst <= x"07DC0080";
end if;
if pc = 30408 then
	inst <= x"820076E8";
end if;
if pc = 30412 then
	inst <= x"0220FFFF";
end if;
if pc = 30416 then
	inst <= x"C17DFFFC";
end if;
if pc = 30420 then
	inst <= x"03DC0080";
end if;
if pc = 30424 then
	inst <= x"037E000C";
end if;
if pc = 30428 then
	inst <= x"C57DFFFC";
end if;
if pc = 30432 then
	inst <= x"8200084C";
end if;
if pc = 30436 then
	inst <= x"07DC0080";
end if;
if pc = 30440 then
	inst <= x"48222000";
end if;
if pc = 30444 then
	inst <= x"C8400044";
end if;
if pc = 30448 then
	inst <= x"48642000";
end if;
if pc = 30452 then
	inst <= x"C03C0000";
end if;
if pc = 30456 then
	inst <= x"CC620000";
end if;
if pc = 30460 then
	inst <= x"C86000A8";
end if;
if pc = 30464 then
	inst <= x"44262000";
end if;
if pc = 30468 then
	inst <= x"48242000";
end if;
if pc = 30472 then
	inst <= x"CC220004";
end if;
if pc = 30476 then
	inst <= x"C1FDFFFC";
end if;
if pc = 30480 then
	inst <= x"C8240000";
end if;
if pc = 30484 then
	inst <= x"C0620014";
end if;
if pc = 30488 then
	inst <= x"C8460000";
end if;
if pc = 30492 then
	inst <= x"44224000";
end if;
if pc = 30496 then
	inst <= x"C8400034";
end if;
if pc = 30500 then
	inst <= x"48624000";
end if;
if pc = 30504 then
	inst <= x"54660000";
end if;
if pc = 30508 then
	inst <= x"8E067748";
end if;
if pc = 30512 then
	inst <= x"58860000";
end if;
if pc = 30516 then
	inst <= x"8A867744";
end if;
if pc = 30520 then
	inst <= x"06660001";
end if;
if pc = 30524 then
	inst <= x"58660000";
end if;
if pc = 30528 then
	inst <= x"82007744";
end if;
if pc = 30532 then
	inst <= x"8200774C";
end if;
if pc = 30536 then
	inst <= x"58660000";
end if;
if pc = 30540 then
	inst <= x"C8800030";
end if;
if pc = 30544 then
	inst <= x"48668000";
end if;
if pc = 30548 then
	inst <= x"44226000";
end if;
if pc = 30552 then
	inst <= x"C860003C";
end if;
if pc = 30556 then
	inst <= x"C8A40008";
end if;
if pc = 30560 then
	inst <= x"C0220014";
end if;
if pc = 30564 then
	inst <= x"C8C20008";
end if;
if pc = 30568 then
	inst <= x"44AAC000";
end if;
if pc = 30572 then
	inst <= x"484A4000";
end if;
if pc = 30576 then
	inst <= x"54240000";
end if;
if pc = 30580 then
	inst <= x"8E047790";
end if;
if pc = 30584 then
	inst <= x"58C20000";
end if;
if pc = 30588 then
	inst <= x"8AC4778C";
end if;
if pc = 30592 then
	inst <= x"06220001";
end if;
if pc = 30596 then
	inst <= x"58420000";
end if;
if pc = 30600 then
	inst <= x"8200778C";
end if;
if pc = 30604 then
	inst <= x"82007794";
end if;
if pc = 30608 then
	inst <= x"58420000";
end if;
if pc = 30612 then
	inst <= x"48448000";
end if;
if pc = 30616 then
	inst <= x"444A4000";
end if;
if pc = 30620 then
	inst <= x"8E2677B4";
end if;
if pc = 30624 then
	inst <= x"8E4677AC";
end if;
if pc = 30628 then
	inst <= x"C8200044";
end if;
if pc = 30632 then
	inst <= x"820077B0";
end if;
if pc = 30636 then
	inst <= x"40200000";
end if;
if pc = 30640 then
	inst <= x"820077C4";
end if;
if pc = 30644 then
	inst <= x"8E4677C0";
end if;
if pc = 30648 then
	inst <= x"40200000";
end if;
if pc = 30652 then
	inst <= x"820077C4";
end if;
if pc = 30656 then
	inst <= x"C8200044";
end if;
if pc = 30660 then
	inst <= x"CC280004";
end if;
if pc = 30664 then
	inst <= x"C1FDFFFC";
end if;
if pc = 30668 then
	inst <= x"8E0277D4";
end if;
if pc = 30672 then
	inst <= x"82007818";
end if;
if pc = 30676 then
	inst <= x"022002EC";
end if;
if pc = 30680 then
	inst <= x"024002D4";
end if;
if pc = 30684 then
	inst <= x"C8820000";
end if;
if pc = 30688 then
	inst <= x"C8A40000";
end if;
if pc = 30692 then
	inst <= x"48A2A000";
end if;
if pc = 30696 then
	inst <= x"4088A000";
end if;
if pc = 30700 then
	inst <= x"CC820000";
end if;
if pc = 30704 then
	inst <= x"C8820004";
end if;
if pc = 30708 then
	inst <= x"C8A40004";
end if;
if pc = 30712 then
	inst <= x"48A2A000";
end if;
if pc = 30716 then
	inst <= x"4088A000";
end if;
if pc = 30720 then
	inst <= x"CC820004";
end if;
if pc = 30724 then
	inst <= x"C8820008";
end if;
if pc = 30728 then
	inst <= x"C8A40008";
end if;
if pc = 30732 then
	inst <= x"4822A000";
end if;
if pc = 30736 then
	inst <= x"40282000";
end if;
if pc = 30740 then
	inst <= x"CC220008";
end if;
if pc = 30744 then
	inst <= x"8E047820";
end if;
if pc = 30748 then
	inst <= x"C1FDFFFC";
end if;
if pc = 30752 then
	inst <= x"48244000";
end if;
if pc = 30756 then
	inst <= x"48222000";
end if;
if pc = 30760 then
	inst <= x"48226000";
end if;
if pc = 30764 then
	inst <= x"022002EC";
end if;
if pc = 30768 then
	inst <= x"C8420000";
end if;
if pc = 30772 then
	inst <= x"40442000";
end if;
if pc = 30776 then
	inst <= x"CC420000";
end if;
if pc = 30780 then
	inst <= x"C8420004";
end if;
if pc = 30784 then
	inst <= x"40442000";
end if;
if pc = 30788 then
	inst <= x"CC420004";
end if;
if pc = 30792 then
	inst <= x"C8420008";
end if;
if pc = 30796 then
	inst <= x"40242000";
end if;
if pc = 30800 then
	inst <= x"CC220008";
end if;
if pc = 30804 then
	inst <= x"C1FDFFFC";
end if;
if pc = 30808 then
	inst <= x"86207A10";
end if;
if pc = 30812 then
	inst <= x"02600370";
end if;
if pc = 30816 then
	inst <= x"22820220";
end if;
if pc = 30820 then
	inst <= x"D0668000";
end if;
if pc = 30824 then
	inst <= x"C0860004";
end if;
if pc = 30828 then
	inst <= x"02A002B4";
end if;
if pc = 30832 then
	inst <= x"C860002C";
end if;
if pc = 30836 then
	inst <= x"CC6A0000";
end if;
if pc = 30840 then
	inst <= x"02C00000";
end if;
if pc = 30844 then
	inst <= x"02E002A8";
end if;
if pc = 30848 then
	inst <= x"C10E0000";
end if;
if pc = 30852 then
	inst <= x"C43C0000";
end if;
if pc = 30856 then
	inst <= x"CC5C0008";
end if;
if pc = 30860 then
	inst <= x"C45C0010";
end if;
if pc = 30864 then
	inst <= x"CC3C0018";
end if;
if pc = 30868 then
	inst <= x"C49C0020";
end if;
if pc = 30872 then
	inst <= x"C4FC0024";
end if;
if pc = 30876 then
	inst <= x"C47C0028";
end if;
if pc = 30880 then
	inst <= x"C4BC002C";
end if;
if pc = 30884 then
	inst <= x"C17DFFFC";
end if;
if pc = 30888 then
	inst <= x"00680000";
end if;
if pc = 30892 then
	inst <= x"00500000";
end if;
if pc = 30896 then
	inst <= x"002C0000";
end if;
if pc = 30900 then
	inst <= x"03DC0038";
end if;
if pc = 30904 then
	inst <= x"037E000C";
end if;
if pc = 30908 then
	inst <= x"C57DFFFC";
end if;
if pc = 30912 then
	inst <= x"820069E8";
end if;
if pc = 30916 then
	inst <= x"07DC0038";
end if;
if pc = 30920 then
	inst <= x"C03C002C";
end if;
if pc = 30924 then
	inst <= x"C8220000";
end if;
if pc = 30928 then
	inst <= x"C8400070";
end if;
if pc = 30932 then
	inst <= x"8E4278E0";
end if;
if pc = 30936 then
	inst <= x"02200000";
end if;
if pc = 30940 then
	inst <= x"820078F4";
end if;
if pc = 30944 then
	inst <= x"C8400028";
end if;
if pc = 30948 then
	inst <= x"8E2478F0";
end if;
if pc = 30952 then
	inst <= x"02200000";
end if;
if pc = 30956 then
	inst <= x"820078F4";
end if;
if pc = 30960 then
	inst <= x"02200001";
end if;
if pc = 30964 then
	inst <= x"822079F8";
end if;
if pc = 30968 then
	inst <= x"022002C4";
end if;
if pc = 30972 then
	inst <= x"C0220000";
end if;
if pc = 30976 then
	inst <= x"22220220";
end if;
if pc = 30980 then
	inst <= x"024002B0";
end if;
if pc = 30984 then
	inst <= x"C0440000";
end if;
if pc = 30988 then
	inst <= x"00224000";
end if;
if pc = 30992 then
	inst <= x"C05C0028";
end if;
if pc = 30996 then
	inst <= x"C0640000";
end if;
if pc = 31000 then
	inst <= x"82267920";
end if;
if pc = 31004 then
	inst <= x"820079F4";
end if;
if pc = 31008 then
	inst <= x"02200000";
end if;
if pc = 31012 then
	inst <= x"C07C0024";
end if;
if pc = 31016 then
	inst <= x"C0660000";
end if;
if pc = 31020 then
	inst <= x"C17DFFFC";
end if;
if pc = 31024 then
	inst <= x"00460000";
end if;
if pc = 31028 then
	inst <= x"03DC0038";
end if;
if pc = 31032 then
	inst <= x"037E000C";
end if;
if pc = 31036 then
	inst <= x"C57DFFFC";
end if;
if pc = 31040 then
	inst <= x"82005414";
end if;
if pc = 31044 then
	inst <= x"07DC0038";
end if;
if pc = 31048 then
	inst <= x"82207950";
end if;
if pc = 31052 then
	inst <= x"820079F4";
end if;
if pc = 31056 then
	inst <= x"022002C8";
end if;
if pc = 31060 then
	inst <= x"C05C0020";
end if;
if pc = 31064 then
	inst <= x"C0640000";
end if;
if pc = 31068 then
	inst <= x"C8220000";
end if;
if pc = 31072 then
	inst <= x"C8460000";
end if;
if pc = 31076 then
	inst <= x"48224000";
end if;
if pc = 31080 then
	inst <= x"C8420004";
end if;
if pc = 31084 then
	inst <= x"C8660004";
end if;
if pc = 31088 then
	inst <= x"48446000";
end if;
if pc = 31092 then
	inst <= x"40224000";
end if;
if pc = 31096 then
	inst <= x"C8420008";
end if;
if pc = 31100 then
	inst <= x"C8660008";
end if;
if pc = 31104 then
	inst <= x"48446000";
end if;
if pc = 31108 then
	inst <= x"40224000";
end if;
if pc = 31112 then
	inst <= x"C03C0028";
end if;
if pc = 31116 then
	inst <= x"C8420008";
end if;
if pc = 31120 then
	inst <= x"C87C0018";
end if;
if pc = 31124 then
	inst <= x"48846000";
end if;
if pc = 31128 then
	inst <= x"48282000";
end if;
if pc = 31132 then
	inst <= x"C0240000";
end if;
if pc = 31136 then
	inst <= x"C05C0010";
end if;
if pc = 31140 then
	inst <= x"C8840000";
end if;
if pc = 31144 then
	inst <= x"C8A20000";
end if;
if pc = 31148 then
	inst <= x"4888A000";
end if;
if pc = 31152 then
	inst <= x"C8A40004";
end if;
if pc = 31156 then
	inst <= x"C8C20004";
end if;
if pc = 31160 then
	inst <= x"48AAC000";
end if;
if pc = 31164 then
	inst <= x"4088A000";
end if;
if pc = 31168 then
	inst <= x"C8A40008";
end if;
if pc = 31172 then
	inst <= x"C8C20008";
end if;
if pc = 31176 then
	inst <= x"48AAC000";
end if;
if pc = 31180 then
	inst <= x"4088A000";
end if;
if pc = 31184 then
	inst <= x"48448000";
end if;
if pc = 31188 then
	inst <= x"C89C0008";
end if;
if pc = 31192 then
	inst <= x"C17DFFFC";
end if;
if pc = 31196 then
	inst <= x"40608000";
end if;
if pc = 31200 then
	inst <= x"03DC0038";
end if;
if pc = 31204 then
	inst <= x"037E000C";
end if;
if pc = 31208 then
	inst <= x"C57DFFFC";
end if;
if pc = 31212 then
	inst <= x"820077CC";
end if;
if pc = 31216 then
	inst <= x"07DC0038";
end if;
if pc = 31220 then
	inst <= x"820079F8";
end if;
if pc = 31224 then
	inst <= x"C03C0000";
end if;
if pc = 31228 then
	inst <= x"06220001";
end if;
if pc = 31232 then
	inst <= x"C83C0018";
end if;
if pc = 31236 then
	inst <= x"C85C0008";
end if;
if pc = 31240 then
	inst <= x"C05C0010";
end if;
if pc = 31244 then
	inst <= x"82007858";
end if;
if pc = 31248 then
	inst <= x"C1FDFFFC";
end if;
if pc = 31252 then
	inst <= x"02800004";
end if;
if pc = 31256 then
	inst <= x"86828030";
end if;
if pc = 31260 then
	inst <= x"C0860008";
end if;
if pc = 31264 then
	inst <= x"02A002B4";
end if;
if pc = 31268 then
	inst <= x"C860002C";
end if;
if pc = 31272 then
	inst <= x"CC6A0000";
end if;
if pc = 31276 then
	inst <= x"02C00000";
end if;
if pc = 31280 then
	inst <= x"02E002A8";
end if;
if pc = 31284 then
	inst <= x"C10E0000";
end if;
if pc = 31288 then
	inst <= x"CC5C0000";
end if;
if pc = 31292 then
	inst <= x"C4FC0008";
end if;
if pc = 31296 then
	inst <= x"C47C000C";
end if;
if pc = 31300 then
	inst <= x"CC3C0010";
end if;
if pc = 31304 then
	inst <= x"C45C0018";
end if;
if pc = 31308 then
	inst <= x"C49C001C";
end if;
if pc = 31312 then
	inst <= x"C43C0020";
end if;
if pc = 31316 then
	inst <= x"C4BC0024";
end if;
if pc = 31320 then
	inst <= x"C17DFFFC";
end if;
if pc = 31324 then
	inst <= x"00640000";
end if;
if pc = 31328 then
	inst <= x"002C0000";
end if;
if pc = 31332 then
	inst <= x"00500000";
end if;
if pc = 31336 then
	inst <= x"03DC0030";
end if;
if pc = 31340 then
	inst <= x"037E000C";
end if;
if pc = 31344 then
	inst <= x"C57DFFFC";
end if;
if pc = 31348 then
	inst <= x"82005E4C";
end if;
if pc = 31352 then
	inst <= x"07DC0030";
end if;
if pc = 31356 then
	inst <= x"C03C0024";
end if;
if pc = 31360 then
	inst <= x"C8220000";
end if;
if pc = 31364 then
	inst <= x"C8400070";
end if;
if pc = 31368 then
	inst <= x"8E427A94";
end if;
if pc = 31372 then
	inst <= x"02400000";
end if;
if pc = 31376 then
	inst <= x"82007AA8";
end if;
if pc = 31380 then
	inst <= x"C8400028";
end if;
if pc = 31384 then
	inst <= x"8E247AA4";
end if;
if pc = 31388 then
	inst <= x"02400000";
end if;
if pc = 31392 then
	inst <= x"82007AA8";
end if;
if pc = 31396 then
	inst <= x"02400001";
end if;
if pc = 31400 then
	inst <= x"82407F8C";
end if;
if pc = 31404 then
	inst <= x"024002C4";
end if;
if pc = 31408 then
	inst <= x"C0440000";
end if;
if pc = 31412 then
	inst <= x"026000C8";
end if;
if pc = 31416 then
	inst <= x"22840220";
end if;
if pc = 31420 then
	inst <= x"D0668000";
end if;
if pc = 31424 then
	inst <= x"C0860008";
end if;
if pc = 31428 then
	inst <= x"C0A6001C";
end if;
if pc = 31432 then
	inst <= x"C82A0000";
end if;
if pc = 31436 then
	inst <= x"C85C0010";
end if;
if pc = 31440 then
	inst <= x"48224000";
end if;
if pc = 31444 then
	inst <= x"C0A60004";
end if;
if pc = 31448 then
	inst <= x"02C00001";
end if;
if pc = 31452 then
	inst <= x"C49C0028";
end if;
if pc = 31456 then
	inst <= x"CC3C0030";
end if;
if pc = 31460 then
	inst <= x"C45C0038";
end if;
if pc = 31464 then
	inst <= x"C47C003C";
end if;
if pc = 31468 then
	inst <= x"82AC7B50";
end if;
if pc = 31472 then
	inst <= x"02C00002";
end if;
if pc = 31476 then
	inst <= x"82AC7B18";
end if;
if pc = 31480 then
	inst <= x"C17DFFFC";
end if;
if pc = 31484 then
	inst <= x"00260000";
end if;
if pc = 31488 then
	inst <= x"03DC0048";
end if;
if pc = 31492 then
	inst <= x"037E000C";
end if;
if pc = 31496 then
	inst <= x"C57DFFFC";
end if;
if pc = 31500 then
	inst <= x"82006F8C";
end if;
if pc = 31504 then
	inst <= x"07DC0048";
end if;
if pc = 31508 then
	inst <= x"82007B4C";
end if;
if pc = 31512 then
	inst <= x"02A002C8";
end if;
if pc = 31516 then
	inst <= x"C0C60010";
end if;
if pc = 31520 then
	inst <= x"C86C0000";
end if;
if pc = 31524 then
	inst <= x"44606000";
end if;
if pc = 31528 then
	inst <= x"CC6A0000";
end if;
if pc = 31532 then
	inst <= x"C0C60010";
end if;
if pc = 31536 then
	inst <= x"C86C0004";
end if;
if pc = 31540 then
	inst <= x"44606000";
end if;
if pc = 31544 then
	inst <= x"CC6A0004";
end if;
if pc = 31548 then
	inst <= x"C0C60010";
end if;
if pc = 31552 then
	inst <= x"C86C0008";
end if;
if pc = 31556 then
	inst <= x"44606000";
end if;
if pc = 31560 then
	inst <= x"CC6A0008";
end if;
if pc = 31564 then
	inst <= x"82007BA4";
end if;
if pc = 31568 then
	inst <= x"02A002B0";
end if;
if pc = 31572 then
	inst <= x"C0AA0000";
end if;
if pc = 31576 then
	inst <= x"02C002C8";
end if;
if pc = 31580 then
	inst <= x"CC0C0000";
end if;
if pc = 31584 then
	inst <= x"CC0C0004";
end if;
if pc = 31588 then
	inst <= x"CC0C0008";
end if;
if pc = 31592 then
	inst <= x"06EA0001";
end if;
if pc = 31596 then
	inst <= x"06AA0001";
end if;
if pc = 31600 then
	inst <= x"22AA0220";
end if;
if pc = 31604 then
	inst <= x"C11C0018";
end if;
if pc = 31608 then
	inst <= x"D870A000";
end if;
if pc = 31612 then
	inst <= x"8A607B94";
end if;
if pc = 31616 then
	inst <= x"8E067B8C";
end if;
if pc = 31620 then
	inst <= x"C860007C";
end if;
if pc = 31624 then
	inst <= x"82007B90";
end if;
if pc = 31628 then
	inst <= x"C86000A8";
end if;
if pc = 31632 then
	inst <= x"82007B98";
end if;
if pc = 31636 then
	inst <= x"40600000";
end if;
if pc = 31640 then
	inst <= x"44606000";
end if;
if pc = 31644 then
	inst <= x"22AE0220";
end if;
if pc = 31648 then
	inst <= x"DC6CA000";
end if;
if pc = 31652 then
	inst <= x"0220030C";
end if;
if pc = 31656 then
	inst <= x"024002B8";
end if;
if pc = 31660 then
	inst <= x"C8240000";
end if;
if pc = 31664 then
	inst <= x"CC220000";
end if;
if pc = 31668 then
	inst <= x"C8240004";
end if;
if pc = 31672 then
	inst <= x"CC220004";
end if;
if pc = 31676 then
	inst <= x"C8240008";
end if;
if pc = 31680 then
	inst <= x"CC220008";
end if;
if pc = 31684 then
	inst <= x"C03C003C";
end if;
if pc = 31688 then
	inst <= x"C45C0040";
end if;
if pc = 31692 then
	inst <= x"C17DFFFC";
end if;
if pc = 31696 then
	inst <= x"03DC004C";
end if;
if pc = 31700 then
	inst <= x"037E000C";
end if;
if pc = 31704 then
	inst <= x"C57DFFFC";
end if;
if pc = 31708 then
	inst <= x"82007158";
end if;
if pc = 31712 then
	inst <= x"07DC004C";
end if;
if pc = 31716 then
	inst <= x"C03C0038";
end if;
if pc = 31720 then
	inst <= x"22220220";
end if;
if pc = 31724 then
	inst <= x"024002B0";
end if;
if pc = 31728 then
	inst <= x"C0440000";
end if;
if pc = 31732 then
	inst <= x"00224000";
end if;
if pc = 31736 then
	inst <= x"C05C0020";
end if;
if pc = 31740 then
	inst <= x"22640220";
end if;
if pc = 31744 then
	inst <= x"C09C001C";
end if;
if pc = 31748 then
	inst <= x"D4286000";
end if;
if pc = 31752 then
	inst <= x"C03C000C";
end if;
if pc = 31756 then
	inst <= x"C0620004";
end if;
if pc = 31760 then
	inst <= x"22A40220";
end if;
if pc = 31764 then
	inst <= x"D066A000";
end if;
if pc = 31768 then
	inst <= x"C0BC0040";
end if;
if pc = 31772 then
	inst <= x"C82A0000";
end if;
if pc = 31776 then
	inst <= x"CC260000";
end if;
if pc = 31780 then
	inst <= x"C82A0004";
end if;
if pc = 31784 then
	inst <= x"CC260004";
end if;
if pc = 31788 then
	inst <= x"C82A0008";
end if;
if pc = 31792 then
	inst <= x"CC260008";
end if;
if pc = 31796 then
	inst <= x"C062000C";
end if;
if pc = 31800 then
	inst <= x"C0DC003C";
end if;
if pc = 31804 then
	inst <= x"C0EC001C";
end if;
if pc = 31808 then
	inst <= x"C82E0000";
end if;
if pc = 31812 then
	inst <= x"C84000A4";
end if;
if pc = 31816 then
	inst <= x"8E247D0C";
end if;
if pc = 31820 then
	inst <= x"02E00001";
end if;
if pc = 31824 then
	inst <= x"23040220";
end if;
if pc = 31828 then
	inst <= x"D4E70000";
end if;
if pc = 31832 then
	inst <= x"C0620010";
end if;
if pc = 31836 then
	inst <= x"22E40220";
end if;
if pc = 31840 then
	inst <= x"D0E6E000";
end if;
if pc = 31844 then
	inst <= x"030002D4";
end if;
if pc = 31848 then
	inst <= x"C8300000";
end if;
if pc = 31852 then
	inst <= x"CC2E0000";
end if;
if pc = 31856 then
	inst <= x"C8300004";
end if;
if pc = 31860 then
	inst <= x"CC2E0004";
end if;
if pc = 31864 then
	inst <= x"C8300008";
end if;
if pc = 31868 then
	inst <= x"CC2E0008";
end if;
if pc = 31872 then
	inst <= x"22E40220";
end if;
if pc = 31876 then
	inst <= x"D066E000";
end if;
if pc = 31880 then
	inst <= x"C8200024";
end if;
if pc = 31884 then
	inst <= x"C47C0044";
end if;
if pc = 31888 then
	inst <= x"C17DFFFC";
end if;
if pc = 31892 then
	inst <= x"03DC0050";
end if;
if pc = 31896 then
	inst <= x"037E000C";
end if;
if pc = 31900 then
	inst <= x"C57DFFFC";
end if;
if pc = 31904 then
	inst <= x"82000844";
end if;
if pc = 31908 then
	inst <= x"07DC0050";
end if;
if pc = 31912 then
	inst <= x"C85C0030";
end if;
if pc = 31916 then
	inst <= x"48224000";
end if;
if pc = 31920 then
	inst <= x"C03C0044";
end if;
if pc = 31924 then
	inst <= x"C8620000";
end if;
if pc = 31928 then
	inst <= x"48662000";
end if;
if pc = 31932 then
	inst <= x"CC620000";
end if;
if pc = 31936 then
	inst <= x"C8620004";
end if;
if pc = 31940 then
	inst <= x"48662000";
end if;
if pc = 31944 then
	inst <= x"CC620004";
end if;
if pc = 31948 then
	inst <= x"C8620008";
end if;
if pc = 31952 then
	inst <= x"48262000";
end if;
if pc = 31956 then
	inst <= x"CC220008";
end if;
if pc = 31960 then
	inst <= x"C03C000C";
end if;
if pc = 31964 then
	inst <= x"C042001C";
end if;
if pc = 31968 then
	inst <= x"C07C0020";
end if;
if pc = 31972 then
	inst <= x"22860220";
end if;
if pc = 31976 then
	inst <= x"D0448000";
end if;
if pc = 31980 then
	inst <= x"028002C8";
end if;
if pc = 31984 then
	inst <= x"C8280000";
end if;
if pc = 31988 then
	inst <= x"CC240000";
end if;
if pc = 31992 then
	inst <= x"C8280004";
end if;
if pc = 31996 then
	inst <= x"CC240004";
end if;
if pc = 32000 then
	inst <= x"C8280008";
end if;
if pc = 32004 then
	inst <= x"CC240008";
end if;
if pc = 32008 then
	inst <= x"82007D18";
end if;
if pc = 32012 then
	inst <= x"02E00000";
end if;
if pc = 32016 then
	inst <= x"23040220";
end if;
if pc = 32020 then
	inst <= x"D4E70000";
end if;
if pc = 32024 then
	inst <= x"C8200020";
end if;
if pc = 32028 then
	inst <= x"024002C8";
end if;
if pc = 32032 then
	inst <= x"C07C0018";
end if;
if pc = 32036 then
	inst <= x"C8460000";
end if;
if pc = 32040 then
	inst <= x"C8640000";
end if;
if pc = 32044 then
	inst <= x"48446000";
end if;
if pc = 32048 then
	inst <= x"C8660004";
end if;
if pc = 32052 then
	inst <= x"C8840004";
end if;
if pc = 32056 then
	inst <= x"48668000";
end if;
if pc = 32060 then
	inst <= x"40446000";
end if;
if pc = 32064 then
	inst <= x"C8660008";
end if;
if pc = 32068 then
	inst <= x"C8840008";
end if;
if pc = 32072 then
	inst <= x"48668000";
end if;
if pc = 32076 then
	inst <= x"40446000";
end if;
if pc = 32080 then
	inst <= x"48224000";
end if;
if pc = 32084 then
	inst <= x"C8460000";
end if;
if pc = 32088 then
	inst <= x"C8640000";
end if;
if pc = 32092 then
	inst <= x"48626000";
end if;
if pc = 32096 then
	inst <= x"40446000";
end if;
if pc = 32100 then
	inst <= x"CC460000";
end if;
if pc = 32104 then
	inst <= x"C8460004";
end if;
if pc = 32108 then
	inst <= x"C8640004";
end if;
if pc = 32112 then
	inst <= x"48626000";
end if;
if pc = 32116 then
	inst <= x"40446000";
end if;
if pc = 32120 then
	inst <= x"CC460004";
end if;
if pc = 32124 then
	inst <= x"C8460008";
end if;
if pc = 32128 then
	inst <= x"C8640008";
end if;
if pc = 32132 then
	inst <= x"48226000";
end if;
if pc = 32136 then
	inst <= x"40242000";
end if;
if pc = 32140 then
	inst <= x"CC260008";
end if;
if pc = 32144 then
	inst <= x"C09C003C";
end if;
if pc = 32148 then
	inst <= x"C0A8001C";
end if;
if pc = 32152 then
	inst <= x"C82A0004";
end if;
if pc = 32156 then
	inst <= x"C85C0010";
end if;
if pc = 32160 then
	inst <= x"48242000";
end if;
if pc = 32164 then
	inst <= x"02A00000";
end if;
if pc = 32168 then
	inst <= x"C0DC0008";
end if;
if pc = 32172 then
	inst <= x"C0CC0000";
end if;
if pc = 32176 then
	inst <= x"CC3C0048";
end if;
if pc = 32180 then
	inst <= x"C45C0050";
end if;
if pc = 32184 then
	inst <= x"C17DFFFC";
end if;
if pc = 32188 then
	inst <= x"004C0000";
end if;
if pc = 32192 then
	inst <= x"002A0000";
end if;
if pc = 32196 then
	inst <= x"03DC005C";
end if;
if pc = 32200 then
	inst <= x"037E000C";
end if;
if pc = 32204 then
	inst <= x"C57DFFFC";
end if;
if pc = 32208 then
	inst <= x"82005414";
end if;
if pc = 32212 then
	inst <= x"07DC005C";
end if;
if pc = 32216 then
	inst <= x"82207DE0";
end if;
if pc = 32220 then
	inst <= x"82007E78";
end if;
if pc = 32224 then
	inst <= x"022001D0";
end if;
if pc = 32228 then
	inst <= x"C05C0050";
end if;
if pc = 32232 then
	inst <= x"C8240000";
end if;
if pc = 32236 then
	inst <= x"C8420000";
end if;
if pc = 32240 then
	inst <= x"48224000";
end if;
if pc = 32244 then
	inst <= x"C8440004";
end if;
if pc = 32248 then
	inst <= x"C8620004";
end if;
if pc = 32252 then
	inst <= x"48446000";
end if;
if pc = 32256 then
	inst <= x"40224000";
end if;
if pc = 32260 then
	inst <= x"C8440008";
end if;
if pc = 32264 then
	inst <= x"C8620008";
end if;
if pc = 32268 then
	inst <= x"48446000";
end if;
if pc = 32272 then
	inst <= x"40224000";
end if;
if pc = 32276 then
	inst <= x"44202000";
end if;
if pc = 32280 then
	inst <= x"C85C0030";
end if;
if pc = 32284 then
	inst <= x"48224000";
end if;
if pc = 32288 then
	inst <= x"C05C0018";
end if;
if pc = 32292 then
	inst <= x"C8640000";
end if;
if pc = 32296 then
	inst <= x"C8820000";
end if;
if pc = 32300 then
	inst <= x"48668000";
end if;
if pc = 32304 then
	inst <= x"C8840004";
end if;
if pc = 32308 then
	inst <= x"C8A20004";
end if;
if pc = 32312 then
	inst <= x"4888A000";
end if;
if pc = 32316 then
	inst <= x"40668000";
end if;
if pc = 32320 then
	inst <= x"C8840008";
end if;
if pc = 32324 then
	inst <= x"C8A20008";
end if;
if pc = 32328 then
	inst <= x"4888A000";
end if;
if pc = 32332 then
	inst <= x"40668000";
end if;
if pc = 32336 then
	inst <= x"44606000";
end if;
if pc = 32340 then
	inst <= x"C89C0048";
end if;
if pc = 32344 then
	inst <= x"C17DFFFC";
end if;
if pc = 32348 then
	inst <= x"40406000";
end if;
if pc = 32352 then
	inst <= x"40608000";
end if;
if pc = 32356 then
	inst <= x"03DC005C";
end if;
if pc = 32360 then
	inst <= x"037E000C";
end if;
if pc = 32364 then
	inst <= x"C57DFFFC";
end if;
if pc = 32368 then
	inst <= x"820077CC";
end if;
if pc = 32372 then
	inst <= x"07DC005C";
end if;
if pc = 32376 then
	inst <= x"02200318";
end if;
if pc = 32380 then
	inst <= x"C05C0040";
end if;
if pc = 32384 then
	inst <= x"C8240000";
end if;
if pc = 32388 then
	inst <= x"CC220000";
end if;
if pc = 32392 then
	inst <= x"C8240004";
end if;
if pc = 32396 then
	inst <= x"CC220004";
end if;
if pc = 32400 then
	inst <= x"C8240008";
end if;
if pc = 32404 then
	inst <= x"CC220008";
end if;
if pc = 32408 then
	inst <= x"022000C4";
end if;
if pc = 32412 then
	inst <= x"C0220000";
end if;
if pc = 32416 then
	inst <= x"06220001";
end if;
if pc = 32420 then
	inst <= x"C17DFFFC";
end if;
if pc = 32424 then
	inst <= x"01240000";
end if;
if pc = 32428 then
	inst <= x"00420000";
end if;
if pc = 32432 then
	inst <= x"00320000";
end if;
if pc = 32436 then
	inst <= x"03DC005C";
end if;
if pc = 32440 then
	inst <= x"037E000C";
end if;
if pc = 32444 then
	inst <= x"C57DFFFC";
end if;
if pc = 32448 then
	inst <= x"8200462C";
end if;
if pc = 32452 then
	inst <= x"07DC005C";
end if;
if pc = 32456 then
	inst <= x"02200640";
end if;
if pc = 32460 then
	inst <= x"C0220000";
end if;
if pc = 32464 then
	inst <= x"06220001";
end if;
if pc = 32468 then
	inst <= x"C83C0030";
end if;
if pc = 32472 then
	inst <= x"C85C0048";
end if;
if pc = 32476 then
	inst <= x"C05C0018";
end if;
if pc = 32480 then
	inst <= x"C17DFFFC";
end if;
if pc = 32484 then
	inst <= x"03DC005C";
end if;
if pc = 32488 then
	inst <= x"037E000C";
end if;
if pc = 32492 then
	inst <= x"C57DFFFC";
end if;
if pc = 32496 then
	inst <= x"82007858";
end if;
if pc = 32500 then
	inst <= x"07DC005C";
end if;
if pc = 32504 then
	inst <= x"C820001C";
end if;
if pc = 32508 then
	inst <= x"C85C0010";
end if;
if pc = 32512 then
	inst <= x"8E247F08";
end if;
if pc = 32516 then
	inst <= x"C1FDFFFC";
end if;
if pc = 32520 then
	inst <= x"02200004";
end if;
if pc = 32524 then
	inst <= x"C05C0020";
end if;
if pc = 32528 then
	inst <= x"86427F18";
end if;
if pc = 32532 then
	inst <= x"82007F2C";
end if;
if pc = 32536 then
	inst <= x"02240001";
end if;
if pc = 32540 then
	inst <= x"0260FFFF";
end if;
if pc = 32544 then
	inst <= x"22220220";
end if;
if pc = 32548 then
	inst <= x"C09C001C";
end if;
if pc = 32552 then
	inst <= x"D4682000";
end if;
if pc = 32556 then
	inst <= x"02200002";
end if;
if pc = 32560 then
	inst <= x"C07C0028";
end if;
if pc = 32564 then
	inst <= x"82627F3C";
end if;
if pc = 32568 then
	inst <= x"82007F88";
end if;
if pc = 32572 then
	inst <= x"C82000A8";
end if;
if pc = 32576 then
	inst <= x"C03C003C";
end if;
if pc = 32580 then
	inst <= x"C022001C";
end if;
if pc = 32584 then
	inst <= x"C8620000";
end if;
if pc = 32588 then
	inst <= x"44226000";
end if;
if pc = 32592 then
	inst <= x"48242000";
end if;
if pc = 32596 then
	inst <= x"02240001";
end if;
if pc = 32600 then
	inst <= x"C05C0024";
end if;
if pc = 32604 then
	inst <= x"C8440000";
end if;
if pc = 32608 then
	inst <= x"C87C0000";
end if;
if pc = 32612 then
	inst <= x"40464000";
end if;
if pc = 32616 then
	inst <= x"C05C0018";
end if;
if pc = 32620 then
	inst <= x"C07C000C";
end if;
if pc = 32624 then
	inst <= x"C17DFFFC";
end if;
if pc = 32628 then
	inst <= x"03DC005C";
end if;
if pc = 32632 then
	inst <= x"037E000C";
end if;
if pc = 32636 then
	inst <= x"C57DFFFC";
end if;
if pc = 32640 then
	inst <= x"82007A14";
end if;
if pc = 32644 then
	inst <= x"07DC005C";
end if;
if pc = 32648 then
	inst <= x"C1FDFFFC";
end if;
if pc = 32652 then
	inst <= x"0220FFFF";
end if;
if pc = 32656 then
	inst <= x"C05C0020";
end if;
if pc = 32660 then
	inst <= x"22640220";
end if;
if pc = 32664 then
	inst <= x"C09C001C";
end if;
if pc = 32668 then
	inst <= x"D4286000";
end if;
if pc = 32672 then
	inst <= x"8240802C";
end if;
if pc = 32676 then
	inst <= x"022001D0";
end if;
if pc = 32680 then
	inst <= x"C05C0018";
end if;
if pc = 32684 then
	inst <= x"C8240000";
end if;
if pc = 32688 then
	inst <= x"C8420000";
end if;
if pc = 32692 then
	inst <= x"48224000";
end if;
if pc = 32696 then
	inst <= x"C8440004";
end if;
if pc = 32700 then
	inst <= x"C8620004";
end if;
if pc = 32704 then
	inst <= x"48446000";
end if;
if pc = 32708 then
	inst <= x"40224000";
end if;
if pc = 32712 then
	inst <= x"C8440008";
end if;
if pc = 32716 then
	inst <= x"C8620008";
end if;
if pc = 32720 then
	inst <= x"48446000";
end if;
if pc = 32724 then
	inst <= x"40224000";
end if;
if pc = 32728 then
	inst <= x"44202000";
end if;
if pc = 32732 then
	inst <= x"8E027FE4";
end if;
if pc = 32736 then
	inst <= x"C1FDFFFC";
end if;
if pc = 32740 then
	inst <= x"48422000";
end if;
if pc = 32744 then
	inst <= x"48242000";
end if;
if pc = 32748 then
	inst <= x"C85C0010";
end if;
if pc = 32752 then
	inst <= x"48224000";
end if;
if pc = 32756 then
	inst <= x"022001DC";
end if;
if pc = 32760 then
	inst <= x"C8420000";
end if;
if pc = 32764 then
	inst <= x"48224000";
end if;
if pc = 32768 then
	inst <= x"022002EC";
end if;
if pc = 32772 then
	inst <= x"C8420000";
end if;
if pc = 32776 then
	inst <= x"40442000";
end if;
if pc = 32780 then
	inst <= x"CC420000";
end if;
if pc = 32784 then
	inst <= x"C8420004";
end if;
if pc = 32788 then
	inst <= x"40442000";
end if;
if pc = 32792 then
	inst <= x"CC420004";
end if;
if pc = 32796 then
	inst <= x"C8420008";
end if;
if pc = 32800 then
	inst <= x"40242000";
end if;
if pc = 32804 then
	inst <= x"CC220008";
end if;
if pc = 32808 then
	inst <= x"C1FDFFFC";
end if;
if pc = 32812 then
	inst <= x"C1FDFFFC";
end if;
if pc = 32816 then
	inst <= x"C1FDFFFC";
end if;
if pc = 32820 then
	inst <= x"024002B4";
end if;
if pc = 32824 then
	inst <= x"C840002C";
end if;
if pc = 32828 then
	inst <= x"CC440000";
end if;
if pc = 32832 then
	inst <= x"02600000";
end if;
if pc = 32836 then
	inst <= x"028002A8";
end if;
if pc = 32840 then
	inst <= x"C0A80000";
end if;
if pc = 32844 then
	inst <= x"CC3C0000";
end if;
if pc = 32848 then
	inst <= x"C49C0008";
end if;
if pc = 32852 then
	inst <= x"C43C000C";
end if;
if pc = 32856 then
	inst <= x"C45C0010";
end if;
if pc = 32860 then
	inst <= x"C17DFFFC";
end if;
if pc = 32864 then
	inst <= x"004A0000";
end if;
if pc = 32868 then
	inst <= x"01260000";
end if;
if pc = 32872 then
	inst <= x"00620000";
end if;
if pc = 32876 then
	inst <= x"00320000";
end if;
if pc = 32880 then
	inst <= x"03DC001C";
end if;
if pc = 32884 then
	inst <= x"037E000C";
end if;
if pc = 32888 then
	inst <= x"C57DFFFC";
end if;
if pc = 32892 then
	inst <= x"820069E8";
end if;
if pc = 32896 then
	inst <= x"07DC001C";
end if;
if pc = 32900 then
	inst <= x"C03C0010";
end if;
if pc = 32904 then
	inst <= x"C8220000";
end if;
if pc = 32908 then
	inst <= x"C8400070";
end if;
if pc = 32912 then
	inst <= x"8E42809C";
end if;
if pc = 32916 then
	inst <= x"02200000";
end if;
if pc = 32920 then
	inst <= x"820080B0";
end if;
if pc = 32924 then
	inst <= x"C8400028";
end if;
if pc = 32928 then
	inst <= x"8E2480AC";
end if;
if pc = 32932 then
	inst <= x"02200000";
end if;
if pc = 32936 then
	inst <= x"820080B0";
end if;
if pc = 32940 then
	inst <= x"02200001";
end if;
if pc = 32944 then
	inst <= x"8220827C";
end if;
if pc = 32948 then
	inst <= x"022000C8";
end if;
if pc = 32952 then
	inst <= x"024002C4";
end if;
if pc = 32956 then
	inst <= x"C0440000";
end if;
if pc = 32960 then
	inst <= x"22440220";
end if;
if pc = 32964 then
	inst <= x"D0224000";
end if;
if pc = 32968 then
	inst <= x"C05C000C";
end if;
if pc = 32972 then
	inst <= x"C0440000";
end if;
if pc = 32976 then
	inst <= x"C0620004";
end if;
if pc = 32980 then
	inst <= x"02800001";
end if;
if pc = 32984 then
	inst <= x"C43C0014";
end if;
if pc = 32988 then
	inst <= x"8268813C";
end if;
if pc = 32992 then
	inst <= x"02400002";
end if;
if pc = 32996 then
	inst <= x"82648104";
end if;
if pc = 33000 then
	inst <= x"C17DFFFC";
end if;
if pc = 33004 then
	inst <= x"03DC0020";
end if;
if pc = 33008 then
	inst <= x"037E000C";
end if;
if pc = 33012 then
	inst <= x"C57DFFFC";
end if;
if pc = 33016 then
	inst <= x"82006F8C";
end if;
if pc = 33020 then
	inst <= x"07DC0020";
end if;
if pc = 33024 then
	inst <= x"82008138";
end if;
if pc = 33028 then
	inst <= x"024002C8";
end if;
if pc = 33032 then
	inst <= x"C0620010";
end if;
if pc = 33036 then
	inst <= x"C8260000";
end if;
if pc = 33040 then
	inst <= x"44202000";
end if;
if pc = 33044 then
	inst <= x"CC240000";
end if;
if pc = 33048 then
	inst <= x"C0620010";
end if;
if pc = 33052 then
	inst <= x"C8260004";
end if;
if pc = 33056 then
	inst <= x"44202000";
end if;
if pc = 33060 then
	inst <= x"CC240004";
end if;
if pc = 33064 then
	inst <= x"C0620010";
end if;
if pc = 33068 then
	inst <= x"C8260008";
end if;
if pc = 33072 then
	inst <= x"44202000";
end if;
if pc = 33076 then
	inst <= x"CC240008";
end if;
if pc = 33080 then
	inst <= x"8200818C";
end if;
if pc = 33084 then
	inst <= x"026002B0";
end if;
if pc = 33088 then
	inst <= x"C0660000";
end if;
if pc = 33092 then
	inst <= x"028002C8";
end if;
if pc = 33096 then
	inst <= x"CC080000";
end if;
if pc = 33100 then
	inst <= x"CC080004";
end if;
if pc = 33104 then
	inst <= x"CC080008";
end if;
if pc = 33108 then
	inst <= x"06A60001";
end if;
if pc = 33112 then
	inst <= x"06660001";
end if;
if pc = 33116 then
	inst <= x"22660220";
end if;
if pc = 33120 then
	inst <= x"D8246000";
end if;
if pc = 33124 then
	inst <= x"8A20817C";
end if;
if pc = 33128 then
	inst <= x"8E028174";
end if;
if pc = 33132 then
	inst <= x"C820007C";
end if;
if pc = 33136 then
	inst <= x"82008178";
end if;
if pc = 33140 then
	inst <= x"C82000A8";
end if;
if pc = 33144 then
	inst <= x"82008180";
end if;
if pc = 33148 then
	inst <= x"40200000";
end if;
if pc = 33152 then
	inst <= x"44202000";
end if;
if pc = 33156 then
	inst <= x"224A0220";
end if;
if pc = 33160 then
	inst <= x"DC284000";
end if;
if pc = 33164 then
	inst <= x"024002B8";
end if;
if pc = 33168 then
	inst <= x"C03C0014";
end if;
if pc = 33172 then
	inst <= x"C17DFFFC";
end if;
if pc = 33176 then
	inst <= x"03DC0020";
end if;
if pc = 33180 then
	inst <= x"037E000C";
end if;
if pc = 33184 then
	inst <= x"C57DFFFC";
end if;
if pc = 33188 then
	inst <= x"82007158";
end if;
if pc = 33192 then
	inst <= x"07DC0020";
end if;
if pc = 33196 then
	inst <= x"02200000";
end if;
if pc = 33200 then
	inst <= x"C05C0008";
end if;
if pc = 33204 then
	inst <= x"C0440000";
end if;
if pc = 33208 then
	inst <= x"C17DFFFC";
end if;
if pc = 33212 then
	inst <= x"03DC0020";
end if;
if pc = 33216 then
	inst <= x"037E000C";
end if;
if pc = 33220 then
	inst <= x"C57DFFFC";
end if;
if pc = 33224 then
	inst <= x"82005414";
end if;
if pc = 33228 then
	inst <= x"07DC0020";
end if;
if pc = 33232 then
	inst <= x"822081D8";
end if;
if pc = 33236 then
	inst <= x"C1FDFFFC";
end if;
if pc = 33240 then
	inst <= x"022002C8";
end if;
if pc = 33244 then
	inst <= x"024001D0";
end if;
if pc = 33248 then
	inst <= x"C8220000";
end if;
if pc = 33252 then
	inst <= x"C8440000";
end if;
if pc = 33256 then
	inst <= x"48224000";
end if;
if pc = 33260 then
	inst <= x"C8420004";
end if;
if pc = 33264 then
	inst <= x"C8640004";
end if;
if pc = 33268 then
	inst <= x"48446000";
end if;
if pc = 33272 then
	inst <= x"40224000";
end if;
if pc = 33276 then
	inst <= x"C8420008";
end if;
if pc = 33280 then
	inst <= x"C8640008";
end if;
if pc = 33284 then
	inst <= x"48446000";
end if;
if pc = 33288 then
	inst <= x"40224000";
end if;
if pc = 33292 then
	inst <= x"44202000";
end if;
if pc = 33296 then
	inst <= x"8E02821C";
end if;
if pc = 33300 then
	inst <= x"40200000";
end if;
if pc = 33304 then
	inst <= x"8200821C";
end if;
if pc = 33308 then
	inst <= x"022002E0";
end if;
if pc = 33312 then
	inst <= x"C85C0000";
end if;
if pc = 33316 then
	inst <= x"48242000";
end if;
if pc = 33320 then
	inst <= x"C05C0014";
end if;
if pc = 33324 then
	inst <= x"C044001C";
end if;
if pc = 33328 then
	inst <= x"C8440000";
end if;
if pc = 33332 then
	inst <= x"48224000";
end if;
if pc = 33336 then
	inst <= x"024002D4";
end if;
if pc = 33340 then
	inst <= x"C8420000";
end if;
if pc = 33344 then
	inst <= x"C8640000";
end if;
if pc = 33348 then
	inst <= x"48626000";
end if;
if pc = 33352 then
	inst <= x"40446000";
end if;
if pc = 33356 then
	inst <= x"CC420000";
end if;
if pc = 33360 then
	inst <= x"C8420004";
end if;
if pc = 33364 then
	inst <= x"C8640004";
end if;
if pc = 33368 then
	inst <= x"48626000";
end if;
if pc = 33372 then
	inst <= x"40446000";
end if;
if pc = 33376 then
	inst <= x"CC420004";
end if;
if pc = 33380 then
	inst <= x"C8420008";
end if;
if pc = 33384 then
	inst <= x"C8640008";
end if;
if pc = 33388 then
	inst <= x"48226000";
end if;
if pc = 33392 then
	inst <= x"40242000";
end if;
if pc = 33396 then
	inst <= x"CC220008";
end if;
if pc = 33400 then
	inst <= x"C1FDFFFC";
end if;
if pc = 33404 then
	inst <= x"C1FDFFFC";
end if;
if pc = 33408 then
	inst <= x"86808490";
end if;
if pc = 33412 then
	inst <= x"22A80220";
end if;
if pc = 33416 then
	inst <= x"D0A2A000";
end if;
if pc = 33420 then
	inst <= x"C0CA0000";
end if;
if pc = 33424 then
	inst <= x"C82C0000";
end if;
if pc = 33428 then
	inst <= x"C8440000";
end if;
if pc = 33432 then
	inst <= x"48224000";
end if;
if pc = 33436 then
	inst <= x"C84C0004";
end if;
if pc = 33440 then
	inst <= x"C8640004";
end if;
if pc = 33444 then
	inst <= x"48446000";
end if;
if pc = 33448 then
	inst <= x"40224000";
end if;
if pc = 33452 then
	inst <= x"C84C0008";
end if;
if pc = 33456 then
	inst <= x"C8640008";
end if;
if pc = 33460 then
	inst <= x"48446000";
end if;
if pc = 33464 then
	inst <= x"40224000";
end if;
if pc = 33468 then
	inst <= x"C47C0000";
end if;
if pc = 33472 then
	inst <= x"C45C0004";
end if;
if pc = 33476 then
	inst <= x"C43C0008";
end if;
if pc = 33480 then
	inst <= x"C49C000C";
end if;
if pc = 33484 then
	inst <= x"8E208320";
end if;
if pc = 33488 then
	inst <= x"C8400018";
end if;
if pc = 33492 then
	inst <= x"C4BC0010";
end if;
if pc = 33496 then
	inst <= x"CC3C0018";
end if;
if pc = 33500 then
	inst <= x"C17DFFFC";
end if;
if pc = 33504 then
	inst <= x"40204000";
end if;
if pc = 33508 then
	inst <= x"03DC0028";
end if;
if pc = 33512 then
	inst <= x"037E000C";
end if;
if pc = 33516 then
	inst <= x"C57DFFFC";
end if;
if pc = 33520 then
	inst <= x"82000844";
end if;
if pc = 33524 then
	inst <= x"07DC0028";
end if;
if pc = 33528 then
	inst <= x"C85C0018";
end if;
if pc = 33532 then
	inst <= x"48242000";
end if;
if pc = 33536 then
	inst <= x"C03C0010";
end if;
if pc = 33540 then
	inst <= x"C17DFFFC";
end if;
if pc = 33544 then
	inst <= x"03DC0028";
end if;
if pc = 33548 then
	inst <= x"037E000C";
end if;
if pc = 33552 then
	inst <= x"C57DFFFC";
end if;
if pc = 33556 then
	inst <= x"82008034";
end if;
if pc = 33560 then
	inst <= x"07DC0028";
end if;
if pc = 33564 then
	inst <= x"82008378";
end if;
if pc = 33568 then
	inst <= x"02A80001";
end if;
if pc = 33572 then
	inst <= x"22AA0220";
end if;
if pc = 33576 then
	inst <= x"D0A2A000";
end if;
if pc = 33580 then
	inst <= x"C8400014";
end if;
if pc = 33584 then
	inst <= x"C4BC0020";
end if;
if pc = 33588 then
	inst <= x"CC3C0018";
end if;
if pc = 33592 then
	inst <= x"C17DFFFC";
end if;
if pc = 33596 then
	inst <= x"40204000";
end if;
if pc = 33600 then
	inst <= x"03DC002C";
end if;
if pc = 33604 then
	inst <= x"037E000C";
end if;
if pc = 33608 then
	inst <= x"C57DFFFC";
end if;
if pc = 33612 then
	inst <= x"82000844";
end if;
if pc = 33616 then
	inst <= x"07DC002C";
end if;
if pc = 33620 then
	inst <= x"C85C0018";
end if;
if pc = 33624 then
	inst <= x"48242000";
end if;
if pc = 33628 then
	inst <= x"C03C0020";
end if;
if pc = 33632 then
	inst <= x"C17DFFFC";
end if;
if pc = 33636 then
	inst <= x"03DC002C";
end if;
if pc = 33640 then
	inst <= x"037E000C";
end if;
if pc = 33644 then
	inst <= x"C57DFFFC";
end if;
if pc = 33648 then
	inst <= x"82008034";
end if;
if pc = 33652 then
	inst <= x"07DC002C";
end if;
if pc = 33656 then
	inst <= x"C03C000C";
end if;
if pc = 33660 then
	inst <= x"06220002";
end if;
if pc = 33664 then
	inst <= x"8620848C";
end if;
if pc = 33668 then
	inst <= x"22420220";
end if;
if pc = 33672 then
	inst <= x"C07C0008";
end if;
if pc = 33676 then
	inst <= x"D0464000";
end if;
if pc = 33680 then
	inst <= x"C0840000";
end if;
if pc = 33684 then
	inst <= x"C8280000";
end if;
if pc = 33688 then
	inst <= x"C0BC0004";
end if;
if pc = 33692 then
	inst <= x"C84A0000";
end if;
if pc = 33696 then
	inst <= x"48224000";
end if;
if pc = 33700 then
	inst <= x"C8480004";
end if;
if pc = 33704 then
	inst <= x"C86A0004";
end if;
if pc = 33708 then
	inst <= x"48446000";
end if;
if pc = 33712 then
	inst <= x"40224000";
end if;
if pc = 33716 then
	inst <= x"C8480008";
end if;
if pc = 33720 then
	inst <= x"C86A0008";
end if;
if pc = 33724 then
	inst <= x"48446000";
end if;
if pc = 33728 then
	inst <= x"40224000";
end if;
if pc = 33732 then
	inst <= x"C43C0024";
end if;
if pc = 33736 then
	inst <= x"8E20841C";
end if;
if pc = 33740 then
	inst <= x"C8400018";
end if;
if pc = 33744 then
	inst <= x"C45C0028";
end if;
if pc = 33748 then
	inst <= x"CC3C0030";
end if;
if pc = 33752 then
	inst <= x"C17DFFFC";
end if;
if pc = 33756 then
	inst <= x"40204000";
end if;
if pc = 33760 then
	inst <= x"03DC0040";
end if;
if pc = 33764 then
	inst <= x"037E000C";
end if;
if pc = 33768 then
	inst <= x"C57DFFFC";
end if;
if pc = 33772 then
	inst <= x"82000844";
end if;
if pc = 33776 then
	inst <= x"07DC0040";
end if;
if pc = 33780 then
	inst <= x"C85C0030";
end if;
if pc = 33784 then
	inst <= x"48242000";
end if;
if pc = 33788 then
	inst <= x"C03C0028";
end if;
if pc = 33792 then
	inst <= x"C17DFFFC";
end if;
if pc = 33796 then
	inst <= x"03DC0040";
end if;
if pc = 33800 then
	inst <= x"037E000C";
end if;
if pc = 33804 then
	inst <= x"C57DFFFC";
end if;
if pc = 33808 then
	inst <= x"82008034";
end if;
if pc = 33812 then
	inst <= x"07DC0040";
end if;
if pc = 33816 then
	inst <= x"82008474";
end if;
if pc = 33820 then
	inst <= x"02420001";
end if;
if pc = 33824 then
	inst <= x"22440220";
end if;
if pc = 33828 then
	inst <= x"D0464000";
end if;
if pc = 33832 then
	inst <= x"C8400014";
end if;
if pc = 33836 then
	inst <= x"C45C0038";
end if;
if pc = 33840 then
	inst <= x"CC3C0030";
end if;
if pc = 33844 then
	inst <= x"C17DFFFC";
end if;
if pc = 33848 then
	inst <= x"40204000";
end if;
if pc = 33852 then
	inst <= x"03DC0044";
end if;
if pc = 33856 then
	inst <= x"037E000C";
end if;
if pc = 33860 then
	inst <= x"C57DFFFC";
end if;
if pc = 33864 then
	inst <= x"82000844";
end if;
if pc = 33868 then
	inst <= x"07DC0044";
end if;
if pc = 33872 then
	inst <= x"C85C0030";
end if;
if pc = 33876 then
	inst <= x"48242000";
end if;
if pc = 33880 then
	inst <= x"C03C0038";
end if;
if pc = 33884 then
	inst <= x"C17DFFFC";
end if;
if pc = 33888 then
	inst <= x"03DC0044";
end if;
if pc = 33892 then
	inst <= x"037E000C";
end if;
if pc = 33896 then
	inst <= x"C57DFFFC";
end if;
if pc = 33900 then
	inst <= x"82008034";
end if;
if pc = 33904 then
	inst <= x"07DC0044";
end if;
if pc = 33908 then
	inst <= x"C03C0024";
end if;
if pc = 33912 then
	inst <= x"06820002";
end if;
if pc = 33916 then
	inst <= x"C03C0008";
end if;
if pc = 33920 then
	inst <= x"C05C0004";
end if;
if pc = 33924 then
	inst <= x"C07C0000";
end if;
if pc = 33928 then
	inst <= x"82008280";
end if;
if pc = 33932 then
	inst <= x"C1FDFFFC";
end if;
if pc = 33936 then
	inst <= x"C1FDFFFC";
end if;
if pc = 33940 then
	inst <= x"C45C0000";
end if;
if pc = 33944 then
	inst <= x"C47C0004";
end if;
if pc = 33948 then
	inst <= x"C43C0008";
end if;
if pc = 33952 then
	inst <= x"82208524";
end if;
if pc = 33956 then
	inst <= x"02800354";
end if;
if pc = 33960 then
	inst <= x"C0880000";
end if;
if pc = 33964 then
	inst <= x"02A00318";
end if;
if pc = 33968 then
	inst <= x"C8260000";
end if;
if pc = 33972 then
	inst <= x"CC2A0000";
end if;
if pc = 33976 then
	inst <= x"C8260004";
end if;
if pc = 33980 then
	inst <= x"CC2A0004";
end if;
if pc = 33984 then
	inst <= x"C8260008";
end if;
if pc = 33988 then
	inst <= x"CC2A0008";
end if;
if pc = 33992 then
	inst <= x"02A000C4";
end if;
if pc = 33996 then
	inst <= x"C0AA0000";
end if;
if pc = 34000 then
	inst <= x"06AA0001";
end if;
if pc = 34004 then
	inst <= x"C49C000C";
end if;
if pc = 34008 then
	inst <= x"C17DFFFC";
end if;
if pc = 34012 then
	inst <= x"004A0000";
end if;
if pc = 34016 then
	inst <= x"00260000";
end if;
if pc = 34020 then
	inst <= x"03DC0018";
end if;
if pc = 34024 then
	inst <= x"037E000C";
end if;
if pc = 34028 then
	inst <= x"C57DFFFC";
end if;
if pc = 34032 then
	inst <= x"8200462C";
end if;
if pc = 34036 then
	inst <= x"07DC0018";
end if;
if pc = 34040 then
	inst <= x"02800076";
end if;
if pc = 34044 then
	inst <= x"C03C000C";
end if;
if pc = 34048 then
	inst <= x"C05C0000";
end if;
if pc = 34052 then
	inst <= x"C07C0004";
end if;
if pc = 34056 then
	inst <= x"C17DFFFC";
end if;
if pc = 34060 then
	inst <= x"03DC0018";
end if;
if pc = 34064 then
	inst <= x"037E000C";
end if;
if pc = 34068 then
	inst <= x"C57DFFFC";
end if;
if pc = 34072 then
	inst <= x"82008280";
end if;
if pc = 34076 then
	inst <= x"07DC0018";
end if;
if pc = 34080 then
	inst <= x"82008524";
end if;
if pc = 34084 then
	inst <= x"02200001";
end if;
if pc = 34088 then
	inst <= x"C05C0008";
end if;
if pc = 34092 then
	inst <= x"824285B4";
end if;
if pc = 34096 then
	inst <= x"02200354";
end if;
if pc = 34100 then
	inst <= x"C0220004";
end if;
if pc = 34104 then
	inst <= x"02600318";
end if;
if pc = 34108 then
	inst <= x"C09C0004";
end if;
if pc = 34112 then
	inst <= x"C8280000";
end if;
if pc = 34116 then
	inst <= x"CC260000";
end if;
if pc = 34120 then
	inst <= x"C8280004";
end if;
if pc = 34124 then
	inst <= x"CC260004";
end if;
if pc = 34128 then
	inst <= x"C8280008";
end if;
if pc = 34132 then
	inst <= x"CC260008";
end if;
if pc = 34136 then
	inst <= x"026000C4";
end if;
if pc = 34140 then
	inst <= x"C0660000";
end if;
if pc = 34144 then
	inst <= x"06660001";
end if;
if pc = 34148 then
	inst <= x"C43C0010";
end if;
if pc = 34152 then
	inst <= x"C17DFFFC";
end if;
if pc = 34156 then
	inst <= x"00460000";
end if;
if pc = 34160 then
	inst <= x"00280000";
end if;
if pc = 34164 then
	inst <= x"03DC001C";
end if;
if pc = 34168 then
	inst <= x"037E000C";
end if;
if pc = 34172 then
	inst <= x"C57DFFFC";
end if;
if pc = 34176 then
	inst <= x"8200462C";
end if;
if pc = 34180 then
	inst <= x"07DC001C";
end if;
if pc = 34184 then
	inst <= x"02800076";
end if;
if pc = 34188 then
	inst <= x"C03C0010";
end if;
if pc = 34192 then
	inst <= x"C05C0000";
end if;
if pc = 34196 then
	inst <= x"C07C0004";
end if;
if pc = 34200 then
	inst <= x"C17DFFFC";
end if;
if pc = 34204 then
	inst <= x"03DC001C";
end if;
if pc = 34208 then
	inst <= x"037E000C";
end if;
if pc = 34212 then
	inst <= x"C57DFFFC";
end if;
if pc = 34216 then
	inst <= x"82008280";
end if;
if pc = 34220 then
	inst <= x"07DC001C";
end if;
if pc = 34224 then
	inst <= x"820085B4";
end if;
if pc = 34228 then
	inst <= x"02200002";
end if;
if pc = 34232 then
	inst <= x"C05C0008";
end if;
if pc = 34236 then
	inst <= x"82428644";
end if;
if pc = 34240 then
	inst <= x"02200354";
end if;
if pc = 34244 then
	inst <= x"C0220008";
end if;
if pc = 34248 then
	inst <= x"02600318";
end if;
if pc = 34252 then
	inst <= x"C09C0004";
end if;
if pc = 34256 then
	inst <= x"C8280000";
end if;
if pc = 34260 then
	inst <= x"CC260000";
end if;
if pc = 34264 then
	inst <= x"C8280004";
end if;
if pc = 34268 then
	inst <= x"CC260004";
end if;
if pc = 34272 then
	inst <= x"C8280008";
end if;
if pc = 34276 then
	inst <= x"CC260008";
end if;
if pc = 34280 then
	inst <= x"026000C4";
end if;
if pc = 34284 then
	inst <= x"C0660000";
end if;
if pc = 34288 then
	inst <= x"06660001";
end if;
if pc = 34292 then
	inst <= x"C43C0014";
end if;
if pc = 34296 then
	inst <= x"C17DFFFC";
end if;
if pc = 34300 then
	inst <= x"00460000";
end if;
if pc = 34304 then
	inst <= x"00280000";
end if;
if pc = 34308 then
	inst <= x"03DC0020";
end if;
if pc = 34312 then
	inst <= x"037E000C";
end if;
if pc = 34316 then
	inst <= x"C57DFFFC";
end if;
if pc = 34320 then
	inst <= x"8200462C";
end if;
if pc = 34324 then
	inst <= x"07DC0020";
end if;
if pc = 34328 then
	inst <= x"02800076";
end if;
if pc = 34332 then
	inst <= x"C03C0014";
end if;
if pc = 34336 then
	inst <= x"C05C0000";
end if;
if pc = 34340 then
	inst <= x"C07C0004";
end if;
if pc = 34344 then
	inst <= x"C17DFFFC";
end if;
if pc = 34348 then
	inst <= x"03DC0020";
end if;
if pc = 34352 then
	inst <= x"037E000C";
end if;
if pc = 34356 then
	inst <= x"C57DFFFC";
end if;
if pc = 34360 then
	inst <= x"82008280";
end if;
if pc = 34364 then
	inst <= x"07DC0020";
end if;
if pc = 34368 then
	inst <= x"82008644";
end if;
if pc = 34372 then
	inst <= x"02200003";
end if;
if pc = 34376 then
	inst <= x"C05C0008";
end if;
if pc = 34380 then
	inst <= x"824286D4";
end if;
if pc = 34384 then
	inst <= x"02200354";
end if;
if pc = 34388 then
	inst <= x"C022000C";
end if;
if pc = 34392 then
	inst <= x"02600318";
end if;
if pc = 34396 then
	inst <= x"C09C0004";
end if;
if pc = 34400 then
	inst <= x"C8280000";
end if;
if pc = 34404 then
	inst <= x"CC260000";
end if;
if pc = 34408 then
	inst <= x"C8280004";
end if;
if pc = 34412 then
	inst <= x"CC260004";
end if;
if pc = 34416 then
	inst <= x"C8280008";
end if;
if pc = 34420 then
	inst <= x"CC260008";
end if;
if pc = 34424 then
	inst <= x"026000C4";
end if;
if pc = 34428 then
	inst <= x"C0660000";
end if;
if pc = 34432 then
	inst <= x"06660001";
end if;
if pc = 34436 then
	inst <= x"C43C0018";
end if;
if pc = 34440 then
	inst <= x"C17DFFFC";
end if;
if pc = 34444 then
	inst <= x"00460000";
end if;
if pc = 34448 then
	inst <= x"00280000";
end if;
if pc = 34452 then
	inst <= x"03DC0024";
end if;
if pc = 34456 then
	inst <= x"037E000C";
end if;
if pc = 34460 then
	inst <= x"C57DFFFC";
end if;
if pc = 34464 then
	inst <= x"8200462C";
end if;
if pc = 34468 then
	inst <= x"07DC0024";
end if;
if pc = 34472 then
	inst <= x"02800076";
end if;
if pc = 34476 then
	inst <= x"C03C0018";
end if;
if pc = 34480 then
	inst <= x"C05C0000";
end if;
if pc = 34484 then
	inst <= x"C07C0004";
end if;
if pc = 34488 then
	inst <= x"C17DFFFC";
end if;
if pc = 34492 then
	inst <= x"03DC0024";
end if;
if pc = 34496 then
	inst <= x"037E000C";
end if;
if pc = 34500 then
	inst <= x"C57DFFFC";
end if;
if pc = 34504 then
	inst <= x"82008280";
end if;
if pc = 34508 then
	inst <= x"07DC0024";
end if;
if pc = 34512 then
	inst <= x"820086D4";
end if;
if pc = 34516 then
	inst <= x"02200004";
end if;
if pc = 34520 then
	inst <= x"C05C0008";
end if;
if pc = 34524 then
	inst <= x"82428748";
end if;
if pc = 34528 then
	inst <= x"02200354";
end if;
if pc = 34532 then
	inst <= x"C0220010";
end if;
if pc = 34536 then
	inst <= x"02400318";
end if;
if pc = 34540 then
	inst <= x"C07C0004";
end if;
if pc = 34544 then
	inst <= x"C8260000";
end if;
if pc = 34548 then
	inst <= x"CC240000";
end if;
if pc = 34552 then
	inst <= x"C8260004";
end if;
if pc = 34556 then
	inst <= x"CC240004";
end if;
if pc = 34560 then
	inst <= x"C8260008";
end if;
if pc = 34564 then
	inst <= x"CC240008";
end if;
if pc = 34568 then
	inst <= x"024000C4";
end if;
if pc = 34572 then
	inst <= x"C0440000";
end if;
if pc = 34576 then
	inst <= x"06440001";
end if;
if pc = 34580 then
	inst <= x"C43C001C";
end if;
if pc = 34584 then
	inst <= x"C17DFFFC";
end if;
if pc = 34588 then
	inst <= x"00260000";
end if;
if pc = 34592 then
	inst <= x"03DC0028";
end if;
if pc = 34596 then
	inst <= x"037E000C";
end if;
if pc = 34600 then
	inst <= x"C57DFFFC";
end if;
if pc = 34604 then
	inst <= x"8200462C";
end if;
if pc = 34608 then
	inst <= x"07DC0028";
end if;
if pc = 34612 then
	inst <= x"02800076";
end if;
if pc = 34616 then
	inst <= x"C03C001C";
end if;
if pc = 34620 then
	inst <= x"C05C0000";
end if;
if pc = 34624 then
	inst <= x"C07C0004";
end if;
if pc = 34628 then
	inst <= x"82008280";
end if;
if pc = 34632 then
	inst <= x"C1FDFFFC";
end if;
if pc = 34636 then
	inst <= x"C0620014";
end if;
if pc = 34640 then
	inst <= x"C082001C";
end if;
if pc = 34644 then
	inst <= x"C0A20004";
end if;
if pc = 34648 then
	inst <= x"C0C20010";
end if;
if pc = 34652 then
	inst <= x"02E002E0";
end if;
if pc = 34656 then
	inst <= x"23040220";
end if;
if pc = 34660 then
	inst <= x"D0670000";
end if;
if pc = 34664 then
	inst <= x"C8260000";
end if;
if pc = 34668 then
	inst <= x"CC2E0000";
end if;
if pc = 34672 then
	inst <= x"C8260004";
end if;
if pc = 34676 then
	inst <= x"CC2E0004";
end if;
if pc = 34680 then
	inst <= x"C8260008";
end if;
if pc = 34684 then
	inst <= x"CC2E0008";
end if;
if pc = 34688 then
	inst <= x"C0220018";
end if;
if pc = 34692 then
	inst <= x"C0220000";
end if;
if pc = 34696 then
	inst <= x"22640220";
end if;
if pc = 34700 then
	inst <= x"D0686000";
end if;
if pc = 34704 then
	inst <= x"22840220";
end if;
if pc = 34708 then
	inst <= x"D08A8000";
end if;
if pc = 34712 then
	inst <= x"C4FC0000";
end if;
if pc = 34716 then
	inst <= x"C4DC0004";
end if;
if pc = 34720 then
	inst <= x"C45C0008";
end if;
if pc = 34724 then
	inst <= x"C47C000C";
end if;
if pc = 34728 then
	inst <= x"C49C0010";
end if;
if pc = 34732 then
	inst <= x"C43C0014";
end if;
if pc = 34736 then
	inst <= x"82208914";
end if;
if pc = 34740 then
	inst <= x"02A00354";
end if;
if pc = 34744 then
	inst <= x"C0AA0000";
end if;
if pc = 34748 then
	inst <= x"03000318";
end if;
if pc = 34752 then
	inst <= x"C8280000";
end if;
if pc = 34756 then
	inst <= x"CC300000";
end if;
if pc = 34760 then
	inst <= x"C8280004";
end if;
if pc = 34764 then
	inst <= x"CC300004";
end if;
if pc = 34768 then
	inst <= x"C8280008";
end if;
if pc = 34772 then
	inst <= x"CC300008";
end if;
if pc = 34776 then
	inst <= x"030000C4";
end if;
if pc = 34780 then
	inst <= x"C1100000";
end if;
if pc = 34784 then
	inst <= x"07100001";
end if;
if pc = 34788 then
	inst <= x"C4BC0018";
end if;
if pc = 34792 then
	inst <= x"C17DFFFC";
end if;
if pc = 34796 then
	inst <= x"00500000";
end if;
if pc = 34800 then
	inst <= x"00280000";
end if;
if pc = 34804 then
	inst <= x"03DC0024";
end if;
if pc = 34808 then
	inst <= x"037E000C";
end if;
if pc = 34812 then
	inst <= x"C57DFFFC";
end if;
if pc = 34816 then
	inst <= x"8200462C";
end if;
if pc = 34820 then
	inst <= x"07DC0024";
end if;
if pc = 34824 then
	inst <= x"C03C0018";
end if;
if pc = 34828 then
	inst <= x"C04201D8";
end if;
if pc = 34832 then
	inst <= x"C0640000";
end if;
if pc = 34836 then
	inst <= x"C8260000";
end if;
if pc = 34840 then
	inst <= x"C09C000C";
end if;
if pc = 34844 then
	inst <= x"C8480000";
end if;
if pc = 34848 then
	inst <= x"48224000";
end if;
if pc = 34852 then
	inst <= x"C8460004";
end if;
if pc = 34856 then
	inst <= x"C8680004";
end if;
if pc = 34860 then
	inst <= x"48446000";
end if;
if pc = 34864 then
	inst <= x"40224000";
end if;
if pc = 34868 then
	inst <= x"C8460008";
end if;
if pc = 34872 then
	inst <= x"C8680008";
end if;
if pc = 34876 then
	inst <= x"48446000";
end if;
if pc = 34880 then
	inst <= x"40224000";
end if;
if pc = 34884 then
	inst <= x"8E208898";
end if;
if pc = 34888 then
	inst <= x"C8400018";
end if;
if pc = 34892 then
	inst <= x"C45C001C";
end if;
if pc = 34896 then
	inst <= x"CC3C0020";
end if;
if pc = 34900 then
	inst <= x"C17DFFFC";
end if;
if pc = 34904 then
	inst <= x"40204000";
end if;
if pc = 34908 then
	inst <= x"03DC0030";
end if;
if pc = 34912 then
	inst <= x"037E000C";
end if;
if pc = 34916 then
	inst <= x"C57DFFFC";
end if;
if pc = 34920 then
	inst <= x"82000844";
end if;
if pc = 34924 then
	inst <= x"07DC0030";
end if;
if pc = 34928 then
	inst <= x"C85C0020";
end if;
if pc = 34932 then
	inst <= x"48242000";
end if;
if pc = 34936 then
	inst <= x"C03C001C";
end if;
if pc = 34940 then
	inst <= x"C17DFFFC";
end if;
if pc = 34944 then
	inst <= x"03DC0030";
end if;
if pc = 34948 then
	inst <= x"037E000C";
end if;
if pc = 34952 then
	inst <= x"C57DFFFC";
end if;
if pc = 34956 then
	inst <= x"82008034";
end if;
if pc = 34960 then
	inst <= x"07DC0030";
end if;
if pc = 34964 then
	inst <= x"820088E8";
end if;
if pc = 34968 then
	inst <= x"C04201DC";
end if;
if pc = 34972 then
	inst <= x"C8400014";
end if;
if pc = 34976 then
	inst <= x"C45C0028";
end if;
if pc = 34980 then
	inst <= x"CC3C0020";
end if;
if pc = 34984 then
	inst <= x"C17DFFFC";
end if;
if pc = 34988 then
	inst <= x"40204000";
end if;
if pc = 34992 then
	inst <= x"03DC0034";
end if;
if pc = 34996 then
	inst <= x"037E000C";
end if;
if pc = 35000 then
	inst <= x"C57DFFFC";
end if;
if pc = 35004 then
	inst <= x"82000844";
end if;
if pc = 35008 then
	inst <= x"07DC0034";
end if;
if pc = 35012 then
	inst <= x"C85C0020";
end if;
if pc = 35016 then
	inst <= x"48242000";
end if;
if pc = 35020 then
	inst <= x"C03C0028";
end if;
if pc = 35024 then
	inst <= x"C17DFFFC";
end if;
if pc = 35028 then
	inst <= x"03DC0034";
end if;
if pc = 35032 then
	inst <= x"037E000C";
end if;
if pc = 35036 then
	inst <= x"C57DFFFC";
end if;
if pc = 35040 then
	inst <= x"82008034";
end if;
if pc = 35044 then
	inst <= x"07DC0034";
end if;
if pc = 35048 then
	inst <= x"02800074";
end if;
if pc = 35052 then
	inst <= x"C03C0018";
end if;
if pc = 35056 then
	inst <= x"C05C000C";
end if;
if pc = 35060 then
	inst <= x"C07C0010";
end if;
if pc = 35064 then
	inst <= x"C17DFFFC";
end if;
if pc = 35068 then
	inst <= x"03DC0034";
end if;
if pc = 35072 then
	inst <= x"037E000C";
end if;
if pc = 35076 then
	inst <= x"C57DFFFC";
end if;
if pc = 35080 then
	inst <= x"82008280";
end if;
if pc = 35084 then
	inst <= x"07DC0034";
end if;
if pc = 35088 then
	inst <= x"82008914";
end if;
if pc = 35092 then
	inst <= x"02200001";
end if;
if pc = 35096 then
	inst <= x"C05C0014";
end if;
if pc = 35100 then
	inst <= x"82428A84";
end if;
if pc = 35104 then
	inst <= x"02200354";
end if;
if pc = 35108 then
	inst <= x"C0220004";
end if;
if pc = 35112 then
	inst <= x"02600318";
end if;
if pc = 35116 then
	inst <= x"C09C0010";
end if;
if pc = 35120 then
	inst <= x"C8280000";
end if;
if pc = 35124 then
	inst <= x"CC260000";
end if;
if pc = 35128 then
	inst <= x"C8280004";
end if;
if pc = 35132 then
	inst <= x"CC260004";
end if;
if pc = 35136 then
	inst <= x"C8280008";
end if;
if pc = 35140 then
	inst <= x"CC260008";
end if;
if pc = 35144 then
	inst <= x"026000C4";
end if;
if pc = 35148 then
	inst <= x"C0660000";
end if;
if pc = 35152 then
	inst <= x"06660001";
end if;
if pc = 35156 then
	inst <= x"C43C002C";
end if;
if pc = 35160 then
	inst <= x"C17DFFFC";
end if;
if pc = 35164 then
	inst <= x"00460000";
end if;
if pc = 35168 then
	inst <= x"00280000";
end if;
if pc = 35172 then
	inst <= x"03DC0038";
end if;
if pc = 35176 then
	inst <= x"037E000C";
end if;
if pc = 35180 then
	inst <= x"C57DFFFC";
end if;
if pc = 35184 then
	inst <= x"8200462C";
end if;
if pc = 35188 then
	inst <= x"07DC0038";
end if;
if pc = 35192 then
	inst <= x"C03C002C";
end if;
if pc = 35196 then
	inst <= x"C04201D8";
end if;
if pc = 35200 then
	inst <= x"C0640000";
end if;
if pc = 35204 then
	inst <= x"C8260000";
end if;
if pc = 35208 then
	inst <= x"C09C000C";
end if;
if pc = 35212 then
	inst <= x"C8480000";
end if;
if pc = 35216 then
	inst <= x"48224000";
end if;
if pc = 35220 then
	inst <= x"C8460004";
end if;
if pc = 35224 then
	inst <= x"C8680004";
end if;
if pc = 35228 then
	inst <= x"48446000";
end if;
if pc = 35232 then
	inst <= x"40224000";
end if;
if pc = 35236 then
	inst <= x"C8460008";
end if;
if pc = 35240 then
	inst <= x"C8680008";
end if;
if pc = 35244 then
	inst <= x"48446000";
end if;
if pc = 35248 then
	inst <= x"40224000";
end if;
if pc = 35252 then
	inst <= x"8E208A08";
end if;
if pc = 35256 then
	inst <= x"C8400018";
end if;
if pc = 35260 then
	inst <= x"C45C0030";
end if;
if pc = 35264 then
	inst <= x"CC3C0038";
end if;
if pc = 35268 then
	inst <= x"C17DFFFC";
end if;
if pc = 35272 then
	inst <= x"40204000";
end if;
if pc = 35276 then
	inst <= x"03DC0048";
end if;
if pc = 35280 then
	inst <= x"037E000C";
end if;
if pc = 35284 then
	inst <= x"C57DFFFC";
end if;
if pc = 35288 then
	inst <= x"82000844";
end if;
if pc = 35292 then
	inst <= x"07DC0048";
end if;
if pc = 35296 then
	inst <= x"C85C0038";
end if;
if pc = 35300 then
	inst <= x"48242000";
end if;
if pc = 35304 then
	inst <= x"C03C0030";
end if;
if pc = 35308 then
	inst <= x"C17DFFFC";
end if;
if pc = 35312 then
	inst <= x"03DC0048";
end if;
if pc = 35316 then
	inst <= x"037E000C";
end if;
if pc = 35320 then
	inst <= x"C57DFFFC";
end if;
if pc = 35324 then
	inst <= x"82008034";
end if;
if pc = 35328 then
	inst <= x"07DC0048";
end if;
if pc = 35332 then
	inst <= x"82008A58";
end if;
if pc = 35336 then
	inst <= x"C04201DC";
end if;
if pc = 35340 then
	inst <= x"C8400014";
end if;
if pc = 35344 then
	inst <= x"C45C0040";
end if;
if pc = 35348 then
	inst <= x"CC3C0038";
end if;
if pc = 35352 then
	inst <= x"C17DFFFC";
end if;
if pc = 35356 then
	inst <= x"40204000";
end if;
if pc = 35360 then
	inst <= x"03DC004C";
end if;
if pc = 35364 then
	inst <= x"037E000C";
end if;
if pc = 35368 then
	inst <= x"C57DFFFC";
end if;
if pc = 35372 then
	inst <= x"82000844";
end if;
if pc = 35376 then
	inst <= x"07DC004C";
end if;
if pc = 35380 then
	inst <= x"C85C0038";
end if;
if pc = 35384 then
	inst <= x"48242000";
end if;
if pc = 35388 then
	inst <= x"C03C0040";
end if;
if pc = 35392 then
	inst <= x"C17DFFFC";
end if;
if pc = 35396 then
	inst <= x"03DC004C";
end if;
if pc = 35400 then
	inst <= x"037E000C";
end if;
if pc = 35404 then
	inst <= x"C57DFFFC";
end if;
if pc = 35408 then
	inst <= x"82008034";
end if;
if pc = 35412 then
	inst <= x"07DC004C";
end if;
if pc = 35416 then
	inst <= x"02800074";
end if;
if pc = 35420 then
	inst <= x"C03C002C";
end if;
if pc = 35424 then
	inst <= x"C05C000C";
end if;
if pc = 35428 then
	inst <= x"C07C0010";
end if;
if pc = 35432 then
	inst <= x"C17DFFFC";
end if;
if pc = 35436 then
	inst <= x"03DC004C";
end if;
if pc = 35440 then
	inst <= x"037E000C";
end if;
if pc = 35444 then
	inst <= x"C57DFFFC";
end if;
if pc = 35448 then
	inst <= x"82008280";
end if;
if pc = 35452 then
	inst <= x"07DC004C";
end if;
if pc = 35456 then
	inst <= x"82008A84";
end if;
if pc = 35460 then
	inst <= x"02200002";
end if;
if pc = 35464 then
	inst <= x"C05C0014";
end if;
if pc = 35468 then
	inst <= x"82428BF4";
end if;
if pc = 35472 then
	inst <= x"02200354";
end if;
if pc = 35476 then
	inst <= x"C0220008";
end if;
if pc = 35480 then
	inst <= x"02600318";
end if;
if pc = 35484 then
	inst <= x"C09C0010";
end if;
if pc = 35488 then
	inst <= x"C8280000";
end if;
if pc = 35492 then
	inst <= x"CC260000";
end if;
if pc = 35496 then
	inst <= x"C8280004";
end if;
if pc = 35500 then
	inst <= x"CC260004";
end if;
if pc = 35504 then
	inst <= x"C8280008";
end if;
if pc = 35508 then
	inst <= x"CC260008";
end if;
if pc = 35512 then
	inst <= x"026000C4";
end if;
if pc = 35516 then
	inst <= x"C0660000";
end if;
if pc = 35520 then
	inst <= x"06660001";
end if;
if pc = 35524 then
	inst <= x"C43C0044";
end if;
if pc = 35528 then
	inst <= x"C17DFFFC";
end if;
if pc = 35532 then
	inst <= x"00460000";
end if;
if pc = 35536 then
	inst <= x"00280000";
end if;
if pc = 35540 then
	inst <= x"03DC0050";
end if;
if pc = 35544 then
	inst <= x"037E000C";
end if;
if pc = 35548 then
	inst <= x"C57DFFFC";
end if;
if pc = 35552 then
	inst <= x"8200462C";
end if;
if pc = 35556 then
	inst <= x"07DC0050";
end if;
if pc = 35560 then
	inst <= x"C03C0044";
end if;
if pc = 35564 then
	inst <= x"C04201D8";
end if;
if pc = 35568 then
	inst <= x"C0640000";
end if;
if pc = 35572 then
	inst <= x"C8260000";
end if;
if pc = 35576 then
	inst <= x"C09C000C";
end if;
if pc = 35580 then
	inst <= x"C8480000";
end if;
if pc = 35584 then
	inst <= x"48224000";
end if;
if pc = 35588 then
	inst <= x"C8460004";
end if;
if pc = 35592 then
	inst <= x"C8680004";
end if;
if pc = 35596 then
	inst <= x"48446000";
end if;
if pc = 35600 then
	inst <= x"40224000";
end if;
if pc = 35604 then
	inst <= x"C8460008";
end if;
if pc = 35608 then
	inst <= x"C8680008";
end if;
if pc = 35612 then
	inst <= x"48446000";
end if;
if pc = 35616 then
	inst <= x"40224000";
end if;
if pc = 35620 then
	inst <= x"8E208B78";
end if;
if pc = 35624 then
	inst <= x"C8400018";
end if;
if pc = 35628 then
	inst <= x"C45C0048";
end if;
if pc = 35632 then
	inst <= x"CC3C0050";
end if;
if pc = 35636 then
	inst <= x"C17DFFFC";
end if;
if pc = 35640 then
	inst <= x"40204000";
end if;
if pc = 35644 then
	inst <= x"03DC0060";
end if;
if pc = 35648 then
	inst <= x"037E000C";
end if;
if pc = 35652 then
	inst <= x"C57DFFFC";
end if;
if pc = 35656 then
	inst <= x"82000844";
end if;
if pc = 35660 then
	inst <= x"07DC0060";
end if;
if pc = 35664 then
	inst <= x"C85C0050";
end if;
if pc = 35668 then
	inst <= x"48242000";
end if;
if pc = 35672 then
	inst <= x"C03C0048";
end if;
if pc = 35676 then
	inst <= x"C17DFFFC";
end if;
if pc = 35680 then
	inst <= x"03DC0060";
end if;
if pc = 35684 then
	inst <= x"037E000C";
end if;
if pc = 35688 then
	inst <= x"C57DFFFC";
end if;
if pc = 35692 then
	inst <= x"82008034";
end if;
if pc = 35696 then
	inst <= x"07DC0060";
end if;
if pc = 35700 then
	inst <= x"82008BC8";
end if;
if pc = 35704 then
	inst <= x"C04201DC";
end if;
if pc = 35708 then
	inst <= x"C8400014";
end if;
if pc = 35712 then
	inst <= x"C45C0058";
end if;
if pc = 35716 then
	inst <= x"CC3C0050";
end if;
if pc = 35720 then
	inst <= x"C17DFFFC";
end if;
if pc = 35724 then
	inst <= x"40204000";
end if;
if pc = 35728 then
	inst <= x"03DC0064";
end if;
if pc = 35732 then
	inst <= x"037E000C";
end if;
if pc = 35736 then
	inst <= x"C57DFFFC";
end if;
if pc = 35740 then
	inst <= x"82000844";
end if;
if pc = 35744 then
	inst <= x"07DC0064";
end if;
if pc = 35748 then
	inst <= x"C85C0050";
end if;
if pc = 35752 then
	inst <= x"48242000";
end if;
if pc = 35756 then
	inst <= x"C03C0058";
end if;
if pc = 35760 then
	inst <= x"C17DFFFC";
end if;
if pc = 35764 then
	inst <= x"03DC0064";
end if;
if pc = 35768 then
	inst <= x"037E000C";
end if;
if pc = 35772 then
	inst <= x"C57DFFFC";
end if;
if pc = 35776 then
	inst <= x"82008034";
end if;
if pc = 35780 then
	inst <= x"07DC0064";
end if;
if pc = 35784 then
	inst <= x"02800074";
end if;
if pc = 35788 then
	inst <= x"C03C0044";
end if;
if pc = 35792 then
	inst <= x"C05C000C";
end if;
if pc = 35796 then
	inst <= x"C07C0010";
end if;
if pc = 35800 then
	inst <= x"C17DFFFC";
end if;
if pc = 35804 then
	inst <= x"03DC0064";
end if;
if pc = 35808 then
	inst <= x"037E000C";
end if;
if pc = 35812 then
	inst <= x"C57DFFFC";
end if;
if pc = 35816 then
	inst <= x"82008280";
end if;
if pc = 35820 then
	inst <= x"07DC0064";
end if;
if pc = 35824 then
	inst <= x"82008BF4";
end if;
if pc = 35828 then
	inst <= x"02200003";
end if;
if pc = 35832 then
	inst <= x"C05C0014";
end if;
if pc = 35836 then
	inst <= x"82428D64";
end if;
if pc = 35840 then
	inst <= x"02200354";
end if;
if pc = 35844 then
	inst <= x"C022000C";
end if;
if pc = 35848 then
	inst <= x"02600318";
end if;
if pc = 35852 then
	inst <= x"C09C0010";
end if;
if pc = 35856 then
	inst <= x"C8280000";
end if;
if pc = 35860 then
	inst <= x"CC260000";
end if;
if pc = 35864 then
	inst <= x"C8280004";
end if;
if pc = 35868 then
	inst <= x"CC260004";
end if;
if pc = 35872 then
	inst <= x"C8280008";
end if;
if pc = 35876 then
	inst <= x"CC260008";
end if;
if pc = 35880 then
	inst <= x"026000C4";
end if;
if pc = 35884 then
	inst <= x"C0660000";
end if;
if pc = 35888 then
	inst <= x"06660001";
end if;
if pc = 35892 then
	inst <= x"C43C005C";
end if;
if pc = 35896 then
	inst <= x"C17DFFFC";
end if;
if pc = 35900 then
	inst <= x"00460000";
end if;
if pc = 35904 then
	inst <= x"00280000";
end if;
if pc = 35908 then
	inst <= x"03DC0068";
end if;
if pc = 35912 then
	inst <= x"037E000C";
end if;
if pc = 35916 then
	inst <= x"C57DFFFC";
end if;
if pc = 35920 then
	inst <= x"8200462C";
end if;
if pc = 35924 then
	inst <= x"07DC0068";
end if;
if pc = 35928 then
	inst <= x"C03C005C";
end if;
if pc = 35932 then
	inst <= x"C04201D8";
end if;
if pc = 35936 then
	inst <= x"C0640000";
end if;
if pc = 35940 then
	inst <= x"C8260000";
end if;
if pc = 35944 then
	inst <= x"C09C000C";
end if;
if pc = 35948 then
	inst <= x"C8480000";
end if;
if pc = 35952 then
	inst <= x"48224000";
end if;
if pc = 35956 then
	inst <= x"C8460004";
end if;
if pc = 35960 then
	inst <= x"C8680004";
end if;
if pc = 35964 then
	inst <= x"48446000";
end if;
if pc = 35968 then
	inst <= x"40224000";
end if;
if pc = 35972 then
	inst <= x"C8460008";
end if;
if pc = 35976 then
	inst <= x"C8680008";
end if;
if pc = 35980 then
	inst <= x"48446000";
end if;
if pc = 35984 then
	inst <= x"40224000";
end if;
if pc = 35988 then
	inst <= x"8E208CE8";
end if;
if pc = 35992 then
	inst <= x"C8400018";
end if;
if pc = 35996 then
	inst <= x"C45C0060";
end if;
if pc = 36000 then
	inst <= x"CC3C0068";
end if;
if pc = 36004 then
	inst <= x"C17DFFFC";
end if;
if pc = 36008 then
	inst <= x"40204000";
end if;
if pc = 36012 then
	inst <= x"03DC0078";
end if;
if pc = 36016 then
	inst <= x"037E000C";
end if;
if pc = 36020 then
	inst <= x"C57DFFFC";
end if;
if pc = 36024 then
	inst <= x"82000844";
end if;
if pc = 36028 then
	inst <= x"07DC0078";
end if;
if pc = 36032 then
	inst <= x"C85C0068";
end if;
if pc = 36036 then
	inst <= x"48242000";
end if;
if pc = 36040 then
	inst <= x"C03C0060";
end if;
if pc = 36044 then
	inst <= x"C17DFFFC";
end if;
if pc = 36048 then
	inst <= x"03DC0078";
end if;
if pc = 36052 then
	inst <= x"037E000C";
end if;
if pc = 36056 then
	inst <= x"C57DFFFC";
end if;
if pc = 36060 then
	inst <= x"82008034";
end if;
if pc = 36064 then
	inst <= x"07DC0078";
end if;
if pc = 36068 then
	inst <= x"82008D38";
end if;
if pc = 36072 then
	inst <= x"C04201DC";
end if;
if pc = 36076 then
	inst <= x"C8400014";
end if;
if pc = 36080 then
	inst <= x"C45C0070";
end if;
if pc = 36084 then
	inst <= x"CC3C0068";
end if;
if pc = 36088 then
	inst <= x"C17DFFFC";
end if;
if pc = 36092 then
	inst <= x"40204000";
end if;
if pc = 36096 then
	inst <= x"03DC007C";
end if;
if pc = 36100 then
	inst <= x"037E000C";
end if;
if pc = 36104 then
	inst <= x"C57DFFFC";
end if;
if pc = 36108 then
	inst <= x"82000844";
end if;
if pc = 36112 then
	inst <= x"07DC007C";
end if;
if pc = 36116 then
	inst <= x"C85C0068";
end if;
if pc = 36120 then
	inst <= x"48242000";
end if;
if pc = 36124 then
	inst <= x"C03C0070";
end if;
if pc = 36128 then
	inst <= x"C17DFFFC";
end if;
if pc = 36132 then
	inst <= x"03DC007C";
end if;
if pc = 36136 then
	inst <= x"037E000C";
end if;
if pc = 36140 then
	inst <= x"C57DFFFC";
end if;
if pc = 36144 then
	inst <= x"82008034";
end if;
if pc = 36148 then
	inst <= x"07DC007C";
end if;
if pc = 36152 then
	inst <= x"02800074";
end if;
if pc = 36156 then
	inst <= x"C03C005C";
end if;
if pc = 36160 then
	inst <= x"C05C000C";
end if;
if pc = 36164 then
	inst <= x"C07C0010";
end if;
if pc = 36168 then
	inst <= x"C17DFFFC";
end if;
if pc = 36172 then
	inst <= x"03DC007C";
end if;
if pc = 36176 then
	inst <= x"037E000C";
end if;
if pc = 36180 then
	inst <= x"C57DFFFC";
end if;
if pc = 36184 then
	inst <= x"82008280";
end if;
if pc = 36188 then
	inst <= x"07DC007C";
end if;
if pc = 36192 then
	inst <= x"82008D64";
end if;
if pc = 36196 then
	inst <= x"02200004";
end if;
if pc = 36200 then
	inst <= x"C05C0014";
end if;
if pc = 36204 then
	inst <= x"82428ED0";
end if;
if pc = 36208 then
	inst <= x"02200354";
end if;
if pc = 36212 then
	inst <= x"C0220010";
end if;
if pc = 36216 then
	inst <= x"02400318";
end if;
if pc = 36220 then
	inst <= x"C07C0010";
end if;
if pc = 36224 then
	inst <= x"C8260000";
end if;
if pc = 36228 then
	inst <= x"CC240000";
end if;
if pc = 36232 then
	inst <= x"C8260004";
end if;
if pc = 36236 then
	inst <= x"CC240004";
end if;
if pc = 36240 then
	inst <= x"C8260008";
end if;
if pc = 36244 then
	inst <= x"CC240008";
end if;
if pc = 36248 then
	inst <= x"024000C4";
end if;
if pc = 36252 then
	inst <= x"C0440000";
end if;
if pc = 36256 then
	inst <= x"06440001";
end if;
if pc = 36260 then
	inst <= x"C43C0074";
end if;
if pc = 36264 then
	inst <= x"C17DFFFC";
end if;
if pc = 36268 then
	inst <= x"00260000";
end if;
if pc = 36272 then
	inst <= x"03DC0080";
end if;
if pc = 36276 then
	inst <= x"037E000C";
end if;
if pc = 36280 then
	inst <= x"C57DFFFC";
end if;
if pc = 36284 then
	inst <= x"8200462C";
end if;
if pc = 36288 then
	inst <= x"07DC0080";
end if;
if pc = 36292 then
	inst <= x"C03C0074";
end if;
if pc = 36296 then
	inst <= x"C04201D8";
end if;
if pc = 36300 then
	inst <= x"C0640000";
end if;
if pc = 36304 then
	inst <= x"C8260000";
end if;
if pc = 36308 then
	inst <= x"C09C000C";
end if;
if pc = 36312 then
	inst <= x"C8480000";
end if;
if pc = 36316 then
	inst <= x"48224000";
end if;
if pc = 36320 then
	inst <= x"C8460004";
end if;
if pc = 36324 then
	inst <= x"C8680004";
end if;
if pc = 36328 then
	inst <= x"48446000";
end if;
if pc = 36332 then
	inst <= x"40224000";
end if;
if pc = 36336 then
	inst <= x"C8460008";
end if;
if pc = 36340 then
	inst <= x"C8680008";
end if;
if pc = 36344 then
	inst <= x"48446000";
end if;
if pc = 36348 then
	inst <= x"40224000";
end if;
if pc = 36352 then
	inst <= x"8E208E54";
end if;
if pc = 36356 then
	inst <= x"C8400018";
end if;
if pc = 36360 then
	inst <= x"C45C0078";
end if;
if pc = 36364 then
	inst <= x"CC3C0080";
end if;
if pc = 36368 then
	inst <= x"C17DFFFC";
end if;
if pc = 36372 then
	inst <= x"40204000";
end if;
if pc = 36376 then
	inst <= x"03DC0090";
end if;
if pc = 36380 then
	inst <= x"037E000C";
end if;
if pc = 36384 then
	inst <= x"C57DFFFC";
end if;
if pc = 36388 then
	inst <= x"82000844";
end if;
if pc = 36392 then
	inst <= x"07DC0090";
end if;
if pc = 36396 then
	inst <= x"C85C0080";
end if;
if pc = 36400 then
	inst <= x"48242000";
end if;
if pc = 36404 then
	inst <= x"C03C0078";
end if;
if pc = 36408 then
	inst <= x"C17DFFFC";
end if;
if pc = 36412 then
	inst <= x"03DC0090";
end if;
if pc = 36416 then
	inst <= x"037E000C";
end if;
if pc = 36420 then
	inst <= x"C57DFFFC";
end if;
if pc = 36424 then
	inst <= x"82008034";
end if;
if pc = 36428 then
	inst <= x"07DC0090";
end if;
if pc = 36432 then
	inst <= x"82008EA4";
end if;
if pc = 36436 then
	inst <= x"C04201DC";
end if;
if pc = 36440 then
	inst <= x"C8400014";
end if;
if pc = 36444 then
	inst <= x"C45C0088";
end if;
if pc = 36448 then
	inst <= x"CC3C0080";
end if;
if pc = 36452 then
	inst <= x"C17DFFFC";
end if;
if pc = 36456 then
	inst <= x"40204000";
end if;
if pc = 36460 then
	inst <= x"03DC0094";
end if;
if pc = 36464 then
	inst <= x"037E000C";
end if;
if pc = 36468 then
	inst <= x"C57DFFFC";
end if;
if pc = 36472 then
	inst <= x"82000844";
end if;
if pc = 36476 then
	inst <= x"07DC0094";
end if;
if pc = 36480 then
	inst <= x"C85C0080";
end if;
if pc = 36484 then
	inst <= x"48242000";
end if;
if pc = 36488 then
	inst <= x"C03C0088";
end if;
if pc = 36492 then
	inst <= x"C17DFFFC";
end if;
if pc = 36496 then
	inst <= x"03DC0094";
end if;
if pc = 36500 then
	inst <= x"037E000C";
end if;
if pc = 36504 then
	inst <= x"C57DFFFC";
end if;
if pc = 36508 then
	inst <= x"82008034";
end if;
if pc = 36512 then
	inst <= x"07DC0094";
end if;
if pc = 36516 then
	inst <= x"02800074";
end if;
if pc = 36520 then
	inst <= x"C03C0074";
end if;
if pc = 36524 then
	inst <= x"C05C000C";
end if;
if pc = 36528 then
	inst <= x"C07C0010";
end if;
if pc = 36532 then
	inst <= x"C17DFFFC";
end if;
if pc = 36536 then
	inst <= x"03DC0094";
end if;
if pc = 36540 then
	inst <= x"037E000C";
end if;
if pc = 36544 then
	inst <= x"C57DFFFC";
end if;
if pc = 36548 then
	inst <= x"82008280";
end if;
if pc = 36552 then
	inst <= x"07DC0094";
end if;
if pc = 36556 then
	inst <= x"82008ED0";
end if;
if pc = 36560 then
	inst <= x"022002EC";
end if;
if pc = 36564 then
	inst <= x"C05C0008";
end if;
if pc = 36568 then
	inst <= x"22440220";
end if;
if pc = 36572 then
	inst <= x"C07C0004";
end if;
if pc = 36576 then
	inst <= x"D0464000";
end if;
if pc = 36580 then
	inst <= x"C8220000";
end if;
if pc = 36584 then
	inst <= x"C8440000";
end if;
if pc = 36588 then
	inst <= x"C07C0000";
end if;
if pc = 36592 then
	inst <= x"C8660000";
end if;
if pc = 36596 then
	inst <= x"48446000";
end if;
if pc = 36600 then
	inst <= x"40224000";
end if;
if pc = 36604 then
	inst <= x"CC220000";
end if;
if pc = 36608 then
	inst <= x"C8220004";
end if;
if pc = 36612 then
	inst <= x"C8440004";
end if;
if pc = 36616 then
	inst <= x"C8660004";
end if;
if pc = 36620 then
	inst <= x"48446000";
end if;
if pc = 36624 then
	inst <= x"40224000";
end if;
if pc = 36628 then
	inst <= x"CC220004";
end if;
if pc = 36632 then
	inst <= x"C8220008";
end if;
if pc = 36636 then
	inst <= x"C8440008";
end if;
if pc = 36640 then
	inst <= x"C8660008";
end if;
if pc = 36644 then
	inst <= x"48446000";
end if;
if pc = 36648 then
	inst <= x"40224000";
end if;
if pc = 36652 then
	inst <= x"CC220008";
end if;
if pc = 36656 then
	inst <= x"C1FDFFFC";
end if;
if pc = 36660 then
	inst <= x"22C20220";
end if;
if pc = 36664 then
	inst <= x"D044C000";
end if;
if pc = 36668 then
	inst <= x"C0440014";
end if;
if pc = 36672 then
	inst <= x"06C20001";
end if;
if pc = 36676 then
	inst <= x"22CC0220";
end if;
if pc = 36680 then
	inst <= x"D0C6C000";
end if;
if pc = 36684 then
	inst <= x"C0CC0014";
end if;
if pc = 36688 then
	inst <= x"22E20220";
end if;
if pc = 36692 then
	inst <= x"D0E6E000";
end if;
if pc = 36696 then
	inst <= x"C0EE0014";
end if;
if pc = 36700 then
	inst <= x"03020001";
end if;
if pc = 36704 then
	inst <= x"23100220";
end if;
if pc = 36708 then
	inst <= x"D1070000";
end if;
if pc = 36712 then
	inst <= x"C1100014";
end if;
if pc = 36716 then
	inst <= x"23220220";
end if;
if pc = 36720 then
	inst <= x"D0892000";
end if;
if pc = 36724 then
	inst <= x"C0880014";
end if;
if pc = 36728 then
	inst <= x"032002E0";
end if;
if pc = 36732 then
	inst <= x"234A0220";
end if;
if pc = 36736 then
	inst <= x"D0454000";
end if;
if pc = 36740 then
	inst <= x"C8240000";
end if;
if pc = 36744 then
	inst <= x"CC320000";
end if;
if pc = 36748 then
	inst <= x"C8240004";
end if;
if pc = 36752 then
	inst <= x"CC320004";
end if;
if pc = 36756 then
	inst <= x"C8240008";
end if;
if pc = 36760 then
	inst <= x"CC320008";
end if;
if pc = 36764 then
	inst <= x"224A0220";
end if;
if pc = 36768 then
	inst <= x"D04C4000";
end if;
if pc = 36772 then
	inst <= x"C8320000";
end if;
if pc = 36776 then
	inst <= x"C8440000";
end if;
if pc = 36780 then
	inst <= x"40224000";
end if;
if pc = 36784 then
	inst <= x"CC320000";
end if;
if pc = 36788 then
	inst <= x"C8320004";
end if;
if pc = 36792 then
	inst <= x"C8440004";
end if;
if pc = 36796 then
	inst <= x"40224000";
end if;
if pc = 36800 then
	inst <= x"CC320004";
end if;
if pc = 36804 then
	inst <= x"C8320008";
end if;
if pc = 36808 then
	inst <= x"C8440008";
end if;
if pc = 36812 then
	inst <= x"40224000";
end if;
if pc = 36816 then
	inst <= x"CC320008";
end if;
if pc = 36820 then
	inst <= x"224A0220";
end if;
if pc = 36824 then
	inst <= x"D04E4000";
end if;
if pc = 36828 then
	inst <= x"C8320000";
end if;
if pc = 36832 then
	inst <= x"C8440000";
end if;
if pc = 36836 then
	inst <= x"40224000";
end if;
if pc = 36840 then
	inst <= x"CC320000";
end if;
if pc = 36844 then
	inst <= x"C8320004";
end if;
if pc = 36848 then
	inst <= x"C8440004";
end if;
if pc = 36852 then
	inst <= x"40224000";
end if;
if pc = 36856 then
	inst <= x"CC320004";
end if;
if pc = 36860 then
	inst <= x"C8320008";
end if;
if pc = 36864 then
	inst <= x"C8440008";
end if;
if pc = 36868 then
	inst <= x"40224000";
end if;
if pc = 36872 then
	inst <= x"CC320008";
end if;
if pc = 36876 then
	inst <= x"224A0220";
end if;
if pc = 36880 then
	inst <= x"D0504000";
end if;
if pc = 36884 then
	inst <= x"C8320000";
end if;
if pc = 36888 then
	inst <= x"C8440000";
end if;
if pc = 36892 then
	inst <= x"40224000";
end if;
if pc = 36896 then
	inst <= x"CC320000";
end if;
if pc = 36900 then
	inst <= x"C8320004";
end if;
if pc = 36904 then
	inst <= x"C8440004";
end if;
if pc = 36908 then
	inst <= x"40224000";
end if;
if pc = 36912 then
	inst <= x"CC320004";
end if;
if pc = 36916 then
	inst <= x"C8320008";
end if;
if pc = 36920 then
	inst <= x"C8440008";
end if;
if pc = 36924 then
	inst <= x"40224000";
end if;
if pc = 36928 then
	inst <= x"CC320008";
end if;
if pc = 36932 then
	inst <= x"224A0220";
end if;
if pc = 36936 then
	inst <= x"D0484000";
end if;
if pc = 36940 then
	inst <= x"C8320000";
end if;
if pc = 36944 then
	inst <= x"C8440000";
end if;
if pc = 36948 then
	inst <= x"40224000";
end if;
if pc = 36952 then
	inst <= x"CC320000";
end if;
if pc = 36956 then
	inst <= x"C8320004";
end if;
if pc = 36960 then
	inst <= x"C8440004";
end if;
if pc = 36964 then
	inst <= x"40224000";
end if;
if pc = 36968 then
	inst <= x"CC320004";
end if;
if pc = 36972 then
	inst <= x"C8320008";
end if;
if pc = 36976 then
	inst <= x"C8440008";
end if;
if pc = 36980 then
	inst <= x"40224000";
end if;
if pc = 36984 then
	inst <= x"CC320008";
end if;
if pc = 36988 then
	inst <= x"22220220";
end if;
if pc = 36992 then
	inst <= x"D0262000";
end if;
if pc = 36996 then
	inst <= x"C0220010";
end if;
if pc = 37000 then
	inst <= x"024002EC";
end if;
if pc = 37004 then
	inst <= x"226A0220";
end if;
if pc = 37008 then
	inst <= x"D0226000";
end if;
if pc = 37012 then
	inst <= x"C8240000";
end if;
if pc = 37016 then
	inst <= x"C8420000";
end if;
if pc = 37020 then
	inst <= x"C8720000";
end if;
if pc = 37024 then
	inst <= x"48446000";
end if;
if pc = 37028 then
	inst <= x"40224000";
end if;
if pc = 37032 then
	inst <= x"CC240000";
end if;
if pc = 37036 then
	inst <= x"C8240004";
end if;
if pc = 37040 then
	inst <= x"C8420004";
end if;
if pc = 37044 then
	inst <= x"C8720004";
end if;
if pc = 37048 then
	inst <= x"48446000";
end if;
if pc = 37052 then
	inst <= x"40224000";
end if;
if pc = 37056 then
	inst <= x"CC240004";
end if;
if pc = 37060 then
	inst <= x"C8240008";
end if;
if pc = 37064 then
	inst <= x"C8420008";
end if;
if pc = 37068 then
	inst <= x"C8720008";
end if;
if pc = 37072 then
	inst <= x"48446000";
end if;
if pc = 37076 then
	inst <= x"40224000";
end if;
if pc = 37080 then
	inst <= x"CC240008";
end if;
if pc = 37084 then
	inst <= x"C1FDFFFC";
end if;
if pc = 37088 then
	inst <= x"02600004";
end if;
if pc = 37092 then
	inst <= x"86649258";
end if;
if pc = 37096 then
	inst <= x"C0620008";
end if;
if pc = 37100 then
	inst <= x"22840220";
end if;
if pc = 37104 then
	inst <= x"D0668000";
end if;
if pc = 37108 then
	inst <= x"86609254";
end if;
if pc = 37112 then
	inst <= x"C062000C";
end if;
if pc = 37116 then
	inst <= x"22840220";
end if;
if pc = 37120 then
	inst <= x"D0668000";
end if;
if pc = 37124 then
	inst <= x"C43C0000";
end if;
if pc = 37128 then
	inst <= x"826091EC";
end if;
if pc = 37132 then
	inst <= x"C0620014";
end if;
if pc = 37136 then
	inst <= x"C082001C";
end if;
if pc = 37140 then
	inst <= x"C0A20004";
end if;
if pc = 37144 then
	inst <= x"C0C20010";
end if;
if pc = 37148 then
	inst <= x"02E002E0";
end if;
if pc = 37152 then
	inst <= x"23040220";
end if;
if pc = 37156 then
	inst <= x"D0670000";
end if;
if pc = 37160 then
	inst <= x"C8260000";
end if;
if pc = 37164 then
	inst <= x"CC2E0000";
end if;
if pc = 37168 then
	inst <= x"C8260004";
end if;
if pc = 37172 then
	inst <= x"CC2E0004";
end if;
if pc = 37176 then
	inst <= x"C8260008";
end if;
if pc = 37180 then
	inst <= x"CC2E0008";
end if;
if pc = 37184 then
	inst <= x"C0620018";
end if;
if pc = 37188 then
	inst <= x"C0660000";
end if;
if pc = 37192 then
	inst <= x"23040220";
end if;
if pc = 37196 then
	inst <= x"D0890000";
end if;
if pc = 37200 then
	inst <= x"23040220";
end if;
if pc = 37204 then
	inst <= x"D0AB0000";
end if;
if pc = 37208 then
	inst <= x"C4FC0004";
end if;
if pc = 37212 then
	inst <= x"C4DC0008";
end if;
if pc = 37216 then
	inst <= x"C45C000C";
end if;
if pc = 37220 then
	inst <= x"C17DFFFC";
end if;
if pc = 37224 then
	inst <= x"00480000";
end if;
if pc = 37228 then
	inst <= x"00260000";
end if;
if pc = 37232 then
	inst <= x"006A0000";
end if;
if pc = 37236 then
	inst <= x"03DC0018";
end if;
if pc = 37240 then
	inst <= x"037E000C";
end if;
if pc = 37244 then
	inst <= x"C57DFFFC";
end if;
if pc = 37248 then
	inst <= x"82008494";
end if;
if pc = 37252 then
	inst <= x"07DC0018";
end if;
if pc = 37256 then
	inst <= x"022002EC";
end if;
if pc = 37260 then
	inst <= x"C05C000C";
end if;
if pc = 37264 then
	inst <= x"22640220";
end if;
if pc = 37268 then
	inst <= x"C09C0008";
end if;
if pc = 37272 then
	inst <= x"D0686000";
end if;
if pc = 37276 then
	inst <= x"C8220000";
end if;
if pc = 37280 then
	inst <= x"C8460000";
end if;
if pc = 37284 then
	inst <= x"C09C0004";
end if;
if pc = 37288 then
	inst <= x"C8680000";
end if;
if pc = 37292 then
	inst <= x"48446000";
end if;
if pc = 37296 then
	inst <= x"40224000";
end if;
if pc = 37300 then
	inst <= x"CC220000";
end if;
if pc = 37304 then
	inst <= x"C8220004";
end if;
if pc = 37308 then
	inst <= x"C8460004";
end if;
if pc = 37312 then
	inst <= x"C8680004";
end if;
if pc = 37316 then
	inst <= x"48446000";
end if;
if pc = 37320 then
	inst <= x"40224000";
end if;
if pc = 37324 then
	inst <= x"CC220004";
end if;
if pc = 37328 then
	inst <= x"C8220008";
end if;
if pc = 37332 then
	inst <= x"C8460008";
end if;
if pc = 37336 then
	inst <= x"C8680008";
end if;
if pc = 37340 then
	inst <= x"48446000";
end if;
if pc = 37344 then
	inst <= x"40224000";
end if;
if pc = 37348 then
	inst <= x"CC220008";
end if;
if pc = 37352 then
	inst <= x"820091EC";
end if;
if pc = 37356 then
	inst <= x"02440001";
end if;
if pc = 37360 then
	inst <= x"02200004";
end if;
if pc = 37364 then
	inst <= x"86249250";
end if;
if pc = 37368 then
	inst <= x"C03C0000";
end if;
if pc = 37372 then
	inst <= x"C0620008";
end if;
if pc = 37376 then
	inst <= x"22840220";
end if;
if pc = 37380 then
	inst <= x"D0668000";
end if;
if pc = 37384 then
	inst <= x"8660924C";
end if;
if pc = 37388 then
	inst <= x"C062000C";
end if;
if pc = 37392 then
	inst <= x"22840220";
end if;
if pc = 37396 then
	inst <= x"D0668000";
end if;
if pc = 37400 then
	inst <= x"C45C0010";
end if;
if pc = 37404 then
	inst <= x"8260923C";
end if;
if pc = 37408 then
	inst <= x"C17DFFFC";
end if;
if pc = 37412 then
	inst <= x"03DC001C";
end if;
if pc = 37416 then
	inst <= x"037E000C";
end if;
if pc = 37420 then
	inst <= x"C57DFFFC";
end if;
if pc = 37424 then
	inst <= x"8200874C";
end if;
if pc = 37428 then
	inst <= x"07DC001C";
end if;
if pc = 37432 then
	inst <= x"8200923C";
end if;
if pc = 37436 then
	inst <= x"C03C0010";
end if;
if pc = 37440 then
	inst <= x"02420001";
end if;
if pc = 37444 then
	inst <= x"C03C0000";
end if;
if pc = 37448 then
	inst <= x"820090E0";
end if;
if pc = 37452 then
	inst <= x"C1FDFFFC";
end if;
if pc = 37456 then
	inst <= x"C1FDFFFC";
end if;
if pc = 37460 then
	inst <= x"C1FDFFFC";
end if;
if pc = 37464 then
	inst <= x"C1FDFFFC";
end if;
if pc = 37468 then
	inst <= x"22E20220";
end if;
if pc = 37472 then
	inst <= x"D0E8E000";
end if;
if pc = 37476 then
	inst <= x"03000004";
end if;
if pc = 37480 then
	inst <= x"870C9528";
end if;
if pc = 37484 then
	inst <= x"C10E0008";
end if;
if pc = 37488 then
	inst <= x"232C0220";
end if;
if pc = 37492 then
	inst <= x"D1112000";
end if;
if pc = 37496 then
	inst <= x"87009524";
end if;
if pc = 37500 then
	inst <= x"C10E0008";
end if;
if pc = 37504 then
	inst <= x"232C0220";
end if;
if pc = 37508 then
	inst <= x"D1112000";
end if;
if pc = 37512 then
	inst <= x"23220220";
end if;
if pc = 37516 then
	inst <= x"D1272000";
end if;
if pc = 37520 then
	inst <= x"C1320008";
end if;
if pc = 37524 then
	inst <= x"234C0220";
end if;
if pc = 37528 then
	inst <= x"D1334000";
end if;
if pc = 37532 then
	inst <= x"833092A8";
end if;
if pc = 37536 then
	inst <= x"03000000";
end if;
if pc = 37540 then
	inst <= x"82009314";
end if;
if pc = 37544 then
	inst <= x"23220220";
end if;
if pc = 37548 then
	inst <= x"D12B2000";
end if;
if pc = 37552 then
	inst <= x"C1320008";
end if;
if pc = 37556 then
	inst <= x"234C0220";
end if;
if pc = 37560 then
	inst <= x"D1334000";
end if;
if pc = 37564 then
	inst <= x"833092C8";
end if;
if pc = 37568 then
	inst <= x"03000000";
end if;
if pc = 37572 then
	inst <= x"82009314";
end if;
if pc = 37576 then
	inst <= x"07220001";
end if;
if pc = 37580 then
	inst <= x"23320220";
end if;
if pc = 37584 then
	inst <= x"D1292000";
end if;
if pc = 37588 then
	inst <= x"C1320008";
end if;
if pc = 37592 then
	inst <= x"234C0220";
end if;
if pc = 37596 then
	inst <= x"D1334000";
end if;
if pc = 37600 then
	inst <= x"833092EC";
end if;
if pc = 37604 then
	inst <= x"03000000";
end if;
if pc = 37608 then
	inst <= x"82009314";
end if;
if pc = 37612 then
	inst <= x"03220001";
end if;
if pc = 37616 then
	inst <= x"23320220";
end if;
if pc = 37620 then
	inst <= x"D1292000";
end if;
if pc = 37624 then
	inst <= x"C1320008";
end if;
if pc = 37628 then
	inst <= x"234C0220";
end if;
if pc = 37632 then
	inst <= x"D1334000";
end if;
if pc = 37636 then
	inst <= x"83309310";
end if;
if pc = 37640 then
	inst <= x"03000000";
end if;
if pc = 37644 then
	inst <= x"82009314";
end if;
if pc = 37648 then
	inst <= x"03000001";
end if;
if pc = 37652 then
	inst <= x"830094B8";
end if;
if pc = 37656 then
	inst <= x"C0EE000C";
end if;
if pc = 37660 then
	inst <= x"230C0220";
end if;
if pc = 37664 then
	inst <= x"D0EF0000";
end if;
if pc = 37668 then
	inst <= x"C45C0000";
end if;
if pc = 37672 then
	inst <= x"C4BC0004";
end if;
if pc = 37676 then
	inst <= x"C47C0008";
end if;
if pc = 37680 then
	inst <= x"C49C000C";
end if;
if pc = 37684 then
	inst <= x"C43C0010";
end if;
if pc = 37688 then
	inst <= x"C4DC0014";
end if;
if pc = 37692 then
	inst <= x"82E0936C";
end if;
if pc = 37696 then
	inst <= x"C17DFFFC";
end if;
if pc = 37700 then
	inst <= x"00460000";
end if;
if pc = 37704 then
	inst <= x"00680000";
end if;
if pc = 37708 then
	inst <= x"008A0000";
end if;
if pc = 37712 then
	inst <= x"00AC0000";
end if;
if pc = 37716 then
	inst <= x"03DC0020";
end if;
if pc = 37720 then
	inst <= x"037E000C";
end if;
if pc = 37724 then
	inst <= x"C57DFFFC";
end if;
if pc = 37728 then
	inst <= x"82008F34";
end if;
if pc = 37732 then
	inst <= x"07DC0020";
end if;
if pc = 37736 then
	inst <= x"8200936C";
end if;
if pc = 37740 then
	inst <= x"C03C0014";
end if;
if pc = 37744 then
	inst <= x"02420001";
end if;
if pc = 37748 then
	inst <= x"C03C0010";
end if;
if pc = 37752 then
	inst <= x"22620220";
end if;
if pc = 37756 then
	inst <= x"C09C000C";
end if;
if pc = 37760 then
	inst <= x"D0686000";
end if;
if pc = 37764 then
	inst <= x"02A00004";
end if;
if pc = 37768 then
	inst <= x"86A494B4";
end if;
if pc = 37772 then
	inst <= x"C0A60008";
end if;
if pc = 37776 then
	inst <= x"22C40220";
end if;
if pc = 37780 then
	inst <= x"D0AAC000";
end if;
if pc = 37784 then
	inst <= x"86A094B0";
end if;
if pc = 37788 then
	inst <= x"C0A60008";
end if;
if pc = 37792 then
	inst <= x"22C40220";
end if;
if pc = 37796 then
	inst <= x"D0AAC000";
end if;
if pc = 37800 then
	inst <= x"22C20220";
end if;
if pc = 37804 then
	inst <= x"C0FC0008";
end if;
if pc = 37808 then
	inst <= x"D0CEC000";
end if;
if pc = 37812 then
	inst <= x"C0CC0008";
end if;
if pc = 37816 then
	inst <= x"23040220";
end if;
if pc = 37820 then
	inst <= x"D0CD0000";
end if;
if pc = 37824 then
	inst <= x"82CA93CC";
end if;
if pc = 37828 then
	inst <= x"02A00000";
end if;
if pc = 37832 then
	inst <= x"8200943C";
end if;
if pc = 37836 then
	inst <= x"22C20220";
end if;
if pc = 37840 then
	inst <= x"C11C0004";
end if;
if pc = 37844 then
	inst <= x"D0D0C000";
end if;
if pc = 37848 then
	inst <= x"C0CC0008";
end if;
if pc = 37852 then
	inst <= x"23240220";
end if;
if pc = 37856 then
	inst <= x"D0CD2000";
end if;
if pc = 37860 then
	inst <= x"82CA93F0";
end if;
if pc = 37864 then
	inst <= x"02A00000";
end if;
if pc = 37868 then
	inst <= x"8200943C";
end if;
if pc = 37872 then
	inst <= x"06C20001";
end if;
if pc = 37876 then
	inst <= x"22CC0220";
end if;
if pc = 37880 then
	inst <= x"D0C8C000";
end if;
if pc = 37884 then
	inst <= x"C0CC0008";
end if;
if pc = 37888 then
	inst <= x"23240220";
end if;
if pc = 37892 then
	inst <= x"D0CD2000";
end if;
if pc = 37896 then
	inst <= x"82CA9414";
end if;
if pc = 37900 then
	inst <= x"02A00000";
end if;
if pc = 37904 then
	inst <= x"8200943C";
end if;
if pc = 37908 then
	inst <= x"02C20001";
end if;
if pc = 37912 then
	inst <= x"22CC0220";
end if;
if pc = 37916 then
	inst <= x"D0C8C000";
end if;
if pc = 37920 then
	inst <= x"C0CC0008";
end if;
if pc = 37924 then
	inst <= x"23240220";
end if;
if pc = 37928 then
	inst <= x"D0CD2000";
end if;
if pc = 37932 then
	inst <= x"82CA9438";
end if;
if pc = 37936 then
	inst <= x"02A00000";
end if;
if pc = 37940 then
	inst <= x"8200943C";
end if;
if pc = 37944 then
	inst <= x"02A00001";
end if;
if pc = 37948 then
	inst <= x"82A094A8";
end if;
if pc = 37952 then
	inst <= x"C066000C";
end if;
if pc = 37956 then
	inst <= x"22A40220";
end if;
if pc = 37960 then
	inst <= x"D066A000";
end if;
if pc = 37964 then
	inst <= x"C45C0018";
end if;
if pc = 37968 then
	inst <= x"82609488";
end if;
if pc = 37972 then
	inst <= x"C07C0004";
end if;
if pc = 37976 then
	inst <= x"C17DFFFC";
end if;
if pc = 37980 then
	inst <= x"00A40000";
end if;
if pc = 37984 then
	inst <= x"004E0000";
end if;
if pc = 37988 then
	inst <= x"01280000";
end if;
if pc = 37992 then
	inst <= x"00860000";
end if;
if pc = 37996 then
	inst <= x"00720000";
end if;
if pc = 38000 then
	inst <= x"03DC0024";
end if;
if pc = 38004 then
	inst <= x"037E000C";
end if;
if pc = 38008 then
	inst <= x"C57DFFFC";
end if;
if pc = 38012 then
	inst <= x"82008F34";
end if;
if pc = 38016 then
	inst <= x"07DC0024";
end if;
if pc = 38020 then
	inst <= x"82009488";
end if;
if pc = 38024 then
	inst <= x"C03C0018";
end if;
if pc = 38028 then
	inst <= x"02C20001";
end if;
if pc = 38032 then
	inst <= x"C03C0010";
end if;
if pc = 38036 then
	inst <= x"C05C0000";
end if;
if pc = 38040 then
	inst <= x"C07C0008";
end if;
if pc = 38044 then
	inst <= x"C09C000C";
end if;
if pc = 38048 then
	inst <= x"C0BC0004";
end if;
if pc = 38052 then
	inst <= x"8200925C";
end if;
if pc = 38056 then
	inst <= x"00260000";
end if;
if pc = 38060 then
	inst <= x"820090E0";
end if;
if pc = 38064 then
	inst <= x"C1FDFFFC";
end if;
if pc = 38068 then
	inst <= x"C1FDFFFC";
end if;
if pc = 38072 then
	inst <= x"02200004";
end if;
if pc = 38076 then
	inst <= x"862C9520";
end if;
if pc = 38080 then
	inst <= x"C02E0008";
end if;
if pc = 38084 then
	inst <= x"224C0220";
end if;
if pc = 38088 then
	inst <= x"D0224000";
end if;
if pc = 38092 then
	inst <= x"8620951C";
end if;
if pc = 38096 then
	inst <= x"C02E000C";
end if;
if pc = 38100 then
	inst <= x"224C0220";
end if;
if pc = 38104 then
	inst <= x"D0224000";
end if;
if pc = 38108 then
	inst <= x"C4FC001C";
end if;
if pc = 38112 then
	inst <= x"C4DC0014";
end if;
if pc = 38116 then
	inst <= x"8220950C";
end if;
if pc = 38120 then
	inst <= x"C17DFFFC";
end if;
if pc = 38124 then
	inst <= x"004C0000";
end if;
if pc = 38128 then
	inst <= x"002E0000";
end if;
if pc = 38132 then
	inst <= x"03DC0028";
end if;
if pc = 38136 then
	inst <= x"037E000C";
end if;
if pc = 38140 then
	inst <= x"C57DFFFC";
end if;
if pc = 38144 then
	inst <= x"8200874C";
end if;
if pc = 38148 then
	inst <= x"07DC0028";
end if;
if pc = 38152 then
	inst <= x"8200950C";
end if;
if pc = 38156 then
	inst <= x"C03C0014";
end if;
if pc = 38160 then
	inst <= x"02420001";
end if;
if pc = 38164 then
	inst <= x"C03C001C";
end if;
if pc = 38168 then
	inst <= x"820090E0";
end if;
if pc = 38172 then
	inst <= x"C1FDFFFC";
end if;
if pc = 38176 then
	inst <= x"C1FDFFFC";
end if;
if pc = 38180 then
	inst <= x"C1FDFFFC";
end if;
if pc = 38184 then
	inst <= x"C1FDFFFC";
end if;
if pc = 38188 then
	inst <= x"02600004";
end if;
if pc = 38192 then
	inst <= x"8664986C";
end if;
if pc = 38196 then
	inst <= x"C0620008";
end if;
if pc = 38200 then
	inst <= x"22840220";
end if;
if pc = 38204 then
	inst <= x"D0668000";
end if;
if pc = 38208 then
	inst <= x"86609868";
end if;
if pc = 38212 then
	inst <= x"C062000C";
end if;
if pc = 38216 then
	inst <= x"22840220";
end if;
if pc = 38220 then
	inst <= x"D0668000";
end if;
if pc = 38224 then
	inst <= x"C45C0000";
end if;
if pc = 38228 then
	inst <= x"8260964C";
end if;
if pc = 38232 then
	inst <= x"C0620018";
end if;
if pc = 38236 then
	inst <= x"C0660000";
end if;
if pc = 38240 then
	inst <= x"028002E0";
end if;
if pc = 38244 then
	inst <= x"CC080000";
end if;
if pc = 38248 then
	inst <= x"CC080004";
end if;
if pc = 38252 then
	inst <= x"CC080008";
end if;
if pc = 38256 then
	inst <= x"C0A2001C";
end if;
if pc = 38260 then
	inst <= x"C0C20004";
end if;
if pc = 38264 then
	inst <= x"02E00354";
end if;
if pc = 38268 then
	inst <= x"22660220";
end if;
if pc = 38272 then
	inst <= x"D06E6000";
end if;
if pc = 38276 then
	inst <= x"22E40220";
end if;
if pc = 38280 then
	inst <= x"D0AAE000";
end if;
if pc = 38284 then
	inst <= x"22E40220";
end if;
if pc = 38288 then
	inst <= x"D0CCE000";
end if;
if pc = 38292 then
	inst <= x"02E00318";
end if;
if pc = 38296 then
	inst <= x"C82C0000";
end if;
if pc = 38300 then
	inst <= x"CC2E0000";
end if;
if pc = 38304 then
	inst <= x"C82C0004";
end if;
if pc = 38308 then
	inst <= x"CC2E0004";
end if;
if pc = 38312 then
	inst <= x"C82C0008";
end if;
if pc = 38316 then
	inst <= x"CC2E0008";
end if;
if pc = 38320 then
	inst <= x"02E000C4";
end if;
if pc = 38324 then
	inst <= x"C0EE0000";
end if;
if pc = 38328 then
	inst <= x"06EE0001";
end if;
if pc = 38332 then
	inst <= x"C49C0004";
end if;
if pc = 38336 then
	inst <= x"C43C0008";
end if;
if pc = 38340 then
	inst <= x"C4DC000C";
end if;
if pc = 38344 then
	inst <= x"C4BC0010";
end if;
if pc = 38348 then
	inst <= x"C47C0014";
end if;
if pc = 38352 then
	inst <= x"C17DFFFC";
end if;
if pc = 38356 then
	inst <= x"004E0000";
end if;
if pc = 38360 then
	inst <= x"002C0000";
end if;
if pc = 38364 then
	inst <= x"03DC0020";
end if;
if pc = 38368 then
	inst <= x"037E000C";
end if;
if pc = 38372 then
	inst <= x"C57DFFFC";
end if;
if pc = 38376 then
	inst <= x"8200462C";
end if;
if pc = 38380 then
	inst <= x"07DC0020";
end if;
if pc = 38384 then
	inst <= x"02800076";
end if;
if pc = 38388 then
	inst <= x"C03C0014";
end if;
if pc = 38392 then
	inst <= x"C05C0010";
end if;
if pc = 38396 then
	inst <= x"C07C000C";
end if;
if pc = 38400 then
	inst <= x"C17DFFFC";
end if;
if pc = 38404 then
	inst <= x"03DC0020";
end if;
if pc = 38408 then
	inst <= x"037E000C";
end if;
if pc = 38412 then
	inst <= x"C57DFFFC";
end if;
if pc = 38416 then
	inst <= x"82008280";
end if;
if pc = 38420 then
	inst <= x"07DC0020";
end if;
if pc = 38424 then
	inst <= x"C03C0008";
end if;
if pc = 38428 then
	inst <= x"C0420014";
end if;
if pc = 38432 then
	inst <= x"C07C0000";
end if;
if pc = 38436 then
	inst <= x"22860220";
end if;
if pc = 38440 then
	inst <= x"D0448000";
end if;
if pc = 38444 then
	inst <= x"C09C0004";
end if;
if pc = 38448 then
	inst <= x"C8280000";
end if;
if pc = 38452 then
	inst <= x"CC240000";
end if;
if pc = 38456 then
	inst <= x"C8280004";
end if;
if pc = 38460 then
	inst <= x"CC240004";
end if;
if pc = 38464 then
	inst <= x"C8280008";
end if;
if pc = 38468 then
	inst <= x"CC240008";
end if;
if pc = 38472 then
	inst <= x"8200964C";
end if;
if pc = 38476 then
	inst <= x"C05C0000";
end if;
if pc = 38480 then
	inst <= x"02440001";
end if;
if pc = 38484 then
	inst <= x"02600004";
end if;
if pc = 38488 then
	inst <= x"86649864";
end if;
if pc = 38492 then
	inst <= x"C0620008";
end if;
if pc = 38496 then
	inst <= x"22840220";
end if;
if pc = 38500 then
	inst <= x"D0668000";
end if;
if pc = 38504 then
	inst <= x"86609860";
end if;
if pc = 38508 then
	inst <= x"C062000C";
end if;
if pc = 38512 then
	inst <= x"22840220";
end if;
if pc = 38516 then
	inst <= x"D0668000";
end if;
if pc = 38520 then
	inst <= x"C45C0018";
end if;
if pc = 38524 then
	inst <= x"82609854";
end if;
if pc = 38528 then
	inst <= x"C0620018";
end if;
if pc = 38532 then
	inst <= x"C0660000";
end if;
if pc = 38536 then
	inst <= x"028002E0";
end if;
if pc = 38540 then
	inst <= x"CC080000";
end if;
if pc = 38544 then
	inst <= x"CC080004";
end if;
if pc = 38548 then
	inst <= x"CC080008";
end if;
if pc = 38552 then
	inst <= x"C0A2001C";
end if;
if pc = 38556 then
	inst <= x"C0C20004";
end if;
if pc = 38560 then
	inst <= x"02E00354";
end if;
if pc = 38564 then
	inst <= x"22660220";
end if;
if pc = 38568 then
	inst <= x"D06E6000";
end if;
if pc = 38572 then
	inst <= x"22E40220";
end if;
if pc = 38576 then
	inst <= x"D0AAE000";
end if;
if pc = 38580 then
	inst <= x"22E40220";
end if;
if pc = 38584 then
	inst <= x"D0CCE000";
end if;
if pc = 38588 then
	inst <= x"02E00318";
end if;
if pc = 38592 then
	inst <= x"C82C0000";
end if;
if pc = 38596 then
	inst <= x"CC2E0000";
end if;
if pc = 38600 then
	inst <= x"C82C0004";
end if;
if pc = 38604 then
	inst <= x"CC2E0004";
end if;
if pc = 38608 then
	inst <= x"C82C0008";
end if;
if pc = 38612 then
	inst <= x"CC2E0008";
end if;
if pc = 38616 then
	inst <= x"02E000C4";
end if;
if pc = 38620 then
	inst <= x"C0EE0000";
end if;
if pc = 38624 then
	inst <= x"06EE0001";
end if;
if pc = 38628 then
	inst <= x"C49C001C";
end if;
if pc = 38632 then
	inst <= x"C43C0008";
end if;
if pc = 38636 then
	inst <= x"C4DC0020";
end if;
if pc = 38640 then
	inst <= x"C4BC0024";
end if;
if pc = 38644 then
	inst <= x"C47C0028";
end if;
if pc = 38648 then
	inst <= x"C17DFFFC";
end if;
if pc = 38652 then
	inst <= x"004E0000";
end if;
if pc = 38656 then
	inst <= x"002C0000";
end if;
if pc = 38660 then
	inst <= x"03DC0034";
end if;
if pc = 38664 then
	inst <= x"037E000C";
end if;
if pc = 38668 then
	inst <= x"C57DFFFC";
end if;
if pc = 38672 then
	inst <= x"8200462C";
end if;
if pc = 38676 then
	inst <= x"07DC0034";
end if;
if pc = 38680 then
	inst <= x"C03C0028";
end if;
if pc = 38684 then
	inst <= x"C04201D8";
end if;
if pc = 38688 then
	inst <= x"C0640000";
end if;
if pc = 38692 then
	inst <= x"C8260000";
end if;
if pc = 38696 then
	inst <= x"C09C0024";
end if;
if pc = 38700 then
	inst <= x"C8480000";
end if;
if pc = 38704 then
	inst <= x"48224000";
end if;
if pc = 38708 then
	inst <= x"C8460004";
end if;
if pc = 38712 then
	inst <= x"C8680004";
end if;
if pc = 38716 then
	inst <= x"48446000";
end if;
if pc = 38720 then
	inst <= x"40224000";
end if;
if pc = 38724 then
	inst <= x"C8460008";
end if;
if pc = 38728 then
	inst <= x"C8680008";
end if;
if pc = 38732 then
	inst <= x"48446000";
end if;
if pc = 38736 then
	inst <= x"40224000";
end if;
if pc = 38740 then
	inst <= x"8E2097A8";
end if;
if pc = 38744 then
	inst <= x"C8400018";
end if;
if pc = 38748 then
	inst <= x"C45C002C";
end if;
if pc = 38752 then
	inst <= x"CC3C0030";
end if;
if pc = 38756 then
	inst <= x"C17DFFFC";
end if;
if pc = 38760 then
	inst <= x"40204000";
end if;
if pc = 38764 then
	inst <= x"03DC0040";
end if;
if pc = 38768 then
	inst <= x"037E000C";
end if;
if pc = 38772 then
	inst <= x"C57DFFFC";
end if;
if pc = 38776 then
	inst <= x"82000844";
end if;
if pc = 38780 then
	inst <= x"07DC0040";
end if;
if pc = 38784 then
	inst <= x"C85C0030";
end if;
if pc = 38788 then
	inst <= x"48242000";
end if;
if pc = 38792 then
	inst <= x"C03C002C";
end if;
if pc = 38796 then
	inst <= x"C17DFFFC";
end if;
if pc = 38800 then
	inst <= x"03DC0040";
end if;
if pc = 38804 then
	inst <= x"037E000C";
end if;
if pc = 38808 then
	inst <= x"C57DFFFC";
end if;
if pc = 38812 then
	inst <= x"82008034";
end if;
if pc = 38816 then
	inst <= x"07DC0040";
end if;
if pc = 38820 then
	inst <= x"820097F8";
end if;
if pc = 38824 then
	inst <= x"C04201DC";
end if;
if pc = 38828 then
	inst <= x"C8400014";
end if;
if pc = 38832 then
	inst <= x"C45C0038";
end if;
if pc = 38836 then
	inst <= x"CC3C0030";
end if;
if pc = 38840 then
	inst <= x"C17DFFFC";
end if;
if pc = 38844 then
	inst <= x"40204000";
end if;
if pc = 38848 then
	inst <= x"03DC0044";
end if;
if pc = 38852 then
	inst <= x"037E000C";
end if;
if pc = 38856 then
	inst <= x"C57DFFFC";
end if;
if pc = 38860 then
	inst <= x"82000844";
end if;
if pc = 38864 then
	inst <= x"07DC0044";
end if;
if pc = 38868 then
	inst <= x"C85C0030";
end if;
if pc = 38872 then
	inst <= x"48242000";
end if;
if pc = 38876 then
	inst <= x"C03C0038";
end if;
if pc = 38880 then
	inst <= x"C17DFFFC";
end if;
if pc = 38884 then
	inst <= x"03DC0044";
end if;
if pc = 38888 then
	inst <= x"037E000C";
end if;
if pc = 38892 then
	inst <= x"C57DFFFC";
end if;
if pc = 38896 then
	inst <= x"82008034";
end if;
if pc = 38900 then
	inst <= x"07DC0044";
end if;
if pc = 38904 then
	inst <= x"02800074";
end if;
if pc = 38908 then
	inst <= x"C03C0028";
end if;
if pc = 38912 then
	inst <= x"C05C0024";
end if;
if pc = 38916 then
	inst <= x"C07C0020";
end if;
if pc = 38920 then
	inst <= x"C17DFFFC";
end if;
if pc = 38924 then
	inst <= x"03DC0044";
end if;
if pc = 38928 then
	inst <= x"037E000C";
end if;
if pc = 38932 then
	inst <= x"C57DFFFC";
end if;
if pc = 38936 then
	inst <= x"82008280";
end if;
if pc = 38940 then
	inst <= x"07DC0044";
end if;
if pc = 38944 then
	inst <= x"C03C0008";
end if;
if pc = 38948 then
	inst <= x"C0420014";
end if;
if pc = 38952 then
	inst <= x"C07C0018";
end if;
if pc = 38956 then
	inst <= x"22860220";
end if;
if pc = 38960 then
	inst <= x"D0448000";
end if;
if pc = 38964 then
	inst <= x"C09C001C";
end if;
if pc = 38968 then
	inst <= x"C8280000";
end if;
if pc = 38972 then
	inst <= x"CC240000";
end if;
if pc = 38976 then
	inst <= x"C8280004";
end if;
if pc = 38980 then
	inst <= x"CC240004";
end if;
if pc = 38984 then
	inst <= x"C8280008";
end if;
if pc = 38988 then
	inst <= x"CC240008";
end if;
if pc = 38992 then
	inst <= x"82009854";
end if;
if pc = 38996 then
	inst <= x"C05C0018";
end if;
if pc = 39000 then
	inst <= x"02440001";
end if;
if pc = 39004 then
	inst <= x"8200952C";
end if;
if pc = 39008 then
	inst <= x"C1FDFFFC";
end if;
if pc = 39012 then
	inst <= x"C1FDFFFC";
end if;
if pc = 39016 then
	inst <= x"C1FDFFFC";
end if;
if pc = 39020 then
	inst <= x"C1FDFFFC";
end if;
if pc = 39024 then
	inst <= x"86409C04";
end if;
if pc = 39028 then
	inst <= x"02800308";
end if;
if pc = 39032 then
	inst <= x"C8880000";
end if;
if pc = 39036 then
	inst <= x"02800300";
end if;
if pc = 39040 then
	inst <= x"C0880000";
end if;
if pc = 39044 then
	inst <= x"04848000";
end if;
if pc = 39048 then
	inst <= x"58A80000";
end if;
if pc = 39052 then
	inst <= x"4888A000";
end if;
if pc = 39056 then
	inst <= x"02800348";
end if;
if pc = 39060 then
	inst <= x"02A00324";
end if;
if pc = 39064 then
	inst <= x"C8AA0000";
end if;
if pc = 39068 then
	inst <= x"48A8A000";
end if;
if pc = 39072 then
	inst <= x"40AA2000";
end if;
if pc = 39076 then
	inst <= x"CCA80000";
end if;
if pc = 39080 then
	inst <= x"C8AA0004";
end if;
if pc = 39084 then
	inst <= x"48A8A000";
end if;
if pc = 39088 then
	inst <= x"40AA4000";
end if;
if pc = 39092 then
	inst <= x"CCA80004";
end if;
if pc = 39096 then
	inst <= x"C8AA0008";
end if;
if pc = 39100 then
	inst <= x"4888A000";
end if;
if pc = 39104 then
	inst <= x"40886000";
end if;
if pc = 39108 then
	inst <= x"CC880008";
end if;
if pc = 39112 then
	inst <= x"02A00000";
end if;
if pc = 39116 then
	inst <= x"CC7C0000";
end if;
if pc = 39120 then
	inst <= x"CC5C0008";
end if;
if pc = 39124 then
	inst <= x"CC3C0010";
end if;
if pc = 39128 then
	inst <= x"C47C0018";
end if;
if pc = 39132 then
	inst <= x"C49C001C";
end if;
if pc = 39136 then
	inst <= x"C43C0020";
end if;
if pc = 39140 then
	inst <= x"C45C0024";
end if;
if pc = 39144 then
	inst <= x"C17DFFFC";
end if;
if pc = 39148 then
	inst <= x"004A0000";
end if;
if pc = 39152 then
	inst <= x"00280000";
end if;
if pc = 39156 then
	inst <= x"03DC0030";
end if;
if pc = 39160 then
	inst <= x"037E000C";
end if;
if pc = 39164 then
	inst <= x"C57DFFFC";
end if;
if pc = 39168 then
	inst <= x"8200161C";
end if;
if pc = 39172 then
	inst <= x"07DC0030";
end if;
if pc = 39176 then
	inst <= x"022002EC";
end if;
if pc = 39180 then
	inst <= x"40400000";
end if;
if pc = 39184 then
	inst <= x"CC020000";
end if;
if pc = 39188 then
	inst <= x"CC020004";
end if;
if pc = 39192 then
	inst <= x"CC020008";
end if;
if pc = 39196 then
	inst <= x"0240030C";
end if;
if pc = 39200 then
	inst <= x"026001C4";
end if;
if pc = 39204 then
	inst <= x"C8260000";
end if;
if pc = 39208 then
	inst <= x"CC240000";
end if;
if pc = 39212 then
	inst <= x"C8260004";
end if;
if pc = 39216 then
	inst <= x"CC240004";
end if;
if pc = 39220 then
	inst <= x"C8260008";
end if;
if pc = 39224 then
	inst <= x"CC240008";
end if;
if pc = 39228 then
	inst <= x"02400000";
end if;
if pc = 39232 then
	inst <= x"C82000A8";
end if;
if pc = 39236 then
	inst <= x"C07C0024";
end if;
if pc = 39240 then
	inst <= x"22860220";
end if;
if pc = 39244 then
	inst <= x"C0BC0020";
end if;
if pc = 39248 then
	inst <= x"D08A8000";
end if;
if pc = 39252 then
	inst <= x"C0DC001C";
end if;
if pc = 39256 then
	inst <= x"C43C0028";
end if;
if pc = 39260 then
	inst <= x"C17DFFFC";
end if;
if pc = 39264 then
	inst <= x"00680000";
end if;
if pc = 39268 then
	inst <= x"00240000";
end if;
if pc = 39272 then
	inst <= x"004C0000";
end if;
if pc = 39276 then
	inst <= x"03DC0034";
end if;
if pc = 39280 then
	inst <= x"037E000C";
end if;
if pc = 39284 then
	inst <= x"C57DFFFC";
end if;
if pc = 39288 then
	inst <= x"82007A14";
end if;
if pc = 39292 then
	inst <= x"07DC0034";
end if;
if pc = 39296 then
	inst <= x"C03C0024";
end if;
if pc = 39300 then
	inst <= x"22420220";
end if;
if pc = 39304 then
	inst <= x"C07C0020";
end if;
if pc = 39308 then
	inst <= x"D0464000";
end if;
if pc = 39312 then
	inst <= x"C0440000";
end if;
if pc = 39316 then
	inst <= x"C09C0028";
end if;
if pc = 39320 then
	inst <= x"C8280000";
end if;
if pc = 39324 then
	inst <= x"CC240000";
end if;
if pc = 39328 then
	inst <= x"C8280004";
end if;
if pc = 39332 then
	inst <= x"CC240004";
end if;
if pc = 39336 then
	inst <= x"C8280008";
end if;
if pc = 39340 then
	inst <= x"CC240008";
end if;
if pc = 39344 then
	inst <= x"22420220";
end if;
if pc = 39348 then
	inst <= x"D0464000";
end if;
if pc = 39352 then
	inst <= x"C0440018";
end if;
if pc = 39356 then
	inst <= x"C09C0018";
end if;
if pc = 39360 then
	inst <= x"C4840000";
end if;
if pc = 39364 then
	inst <= x"22420220";
end if;
if pc = 39368 then
	inst <= x"D0464000";
end if;
if pc = 39372 then
	inst <= x"C0A40008";
end if;
if pc = 39376 then
	inst <= x"C0AA0000";
end if;
if pc = 39380 then
	inst <= x"86A09BCC";
end if;
if pc = 39384 then
	inst <= x"C0A4000C";
end if;
if pc = 39388 then
	inst <= x"C0AA0000";
end if;
if pc = 39392 then
	inst <= x"C45C002C";
end if;
if pc = 39396 then
	inst <= x"82A09BA8";
end if;
if pc = 39400 then
	inst <= x"C0A40018";
end if;
if pc = 39404 then
	inst <= x"C0AA0000";
end if;
if pc = 39408 then
	inst <= x"02C002E0";
end if;
if pc = 39412 then
	inst <= x"CC0C0000";
end if;
if pc = 39416 then
	inst <= x"CC0C0004";
end if;
if pc = 39420 then
	inst <= x"CC0C0008";
end if;
if pc = 39424 then
	inst <= x"C0E4001C";
end if;
if pc = 39428 then
	inst <= x"C1040004";
end if;
if pc = 39432 then
	inst <= x"03200354";
end if;
if pc = 39436 then
	inst <= x"22AA0220";
end if;
if pc = 39440 then
	inst <= x"D0B2A000";
end if;
if pc = 39444 then
	inst <= x"C0EE0000";
end if;
if pc = 39448 then
	inst <= x"C1100000";
end if;
if pc = 39452 then
	inst <= x"03200318";
end if;
if pc = 39456 then
	inst <= x"C8300000";
end if;
if pc = 39460 then
	inst <= x"CC320000";
end if;
if pc = 39464 then
	inst <= x"C8300004";
end if;
if pc = 39468 then
	inst <= x"CC320004";
end if;
if pc = 39472 then
	inst <= x"C8300008";
end if;
if pc = 39476 then
	inst <= x"CC320008";
end if;
if pc = 39480 then
	inst <= x"032000C4";
end if;
if pc = 39484 then
	inst <= x"C1320000";
end if;
if pc = 39488 then
	inst <= x"07320001";
end if;
if pc = 39492 then
	inst <= x"C4DC0030";
end if;
if pc = 39496 then
	inst <= x"C51C0034";
end if;
if pc = 39500 then
	inst <= x"C4FC0038";
end if;
if pc = 39504 then
	inst <= x"C4BC003C";
end if;
if pc = 39508 then
	inst <= x"C17DFFFC";
end if;
if pc = 39512 then
	inst <= x"00520000";
end if;
if pc = 39516 then
	inst <= x"00300000";
end if;
if pc = 39520 then
	inst <= x"03DC0048";
end if;
if pc = 39524 then
	inst <= x"037E000C";
end if;
if pc = 39528 then
	inst <= x"C57DFFFC";
end if;
if pc = 39532 then
	inst <= x"8200462C";
end if;
if pc = 39536 then
	inst <= x"07DC0048";
end if;
if pc = 39540 then
	inst <= x"C03C003C";
end if;
if pc = 39544 then
	inst <= x"C04201D8";
end if;
if pc = 39548 then
	inst <= x"C0640000";
end if;
if pc = 39552 then
	inst <= x"C8260000";
end if;
if pc = 39556 then
	inst <= x"C09C0038";
end if;
if pc = 39560 then
	inst <= x"C8480000";
end if;
if pc = 39564 then
	inst <= x"48224000";
end if;
if pc = 39568 then
	inst <= x"C8460004";
end if;
if pc = 39572 then
	inst <= x"C8680004";
end if;
if pc = 39576 then
	inst <= x"48446000";
end if;
if pc = 39580 then
	inst <= x"40224000";
end if;
if pc = 39584 then
	inst <= x"C8460008";
end if;
if pc = 39588 then
	inst <= x"C8680008";
end if;
if pc = 39592 then
	inst <= x"48446000";
end if;
if pc = 39596 then
	inst <= x"40224000";
end if;
if pc = 39600 then
	inst <= x"8E209B04";
end if;
if pc = 39604 then
	inst <= x"C8400018";
end if;
if pc = 39608 then
	inst <= x"C45C0040";
end if;
if pc = 39612 then
	inst <= x"CC3C0048";
end if;
if pc = 39616 then
	inst <= x"C17DFFFC";
end if;
if pc = 39620 then
	inst <= x"40204000";
end if;
if pc = 39624 then
	inst <= x"03DC0058";
end if;
if pc = 39628 then
	inst <= x"037E000C";
end if;
if pc = 39632 then
	inst <= x"C57DFFFC";
end if;
if pc = 39636 then
	inst <= x"82000844";
end if;
if pc = 39640 then
	inst <= x"07DC0058";
end if;
if pc = 39644 then
	inst <= x"C85C0048";
end if;
if pc = 39648 then
	inst <= x"48242000";
end if;
if pc = 39652 then
	inst <= x"C03C0040";
end if;
if pc = 39656 then
	inst <= x"C17DFFFC";
end if;
if pc = 39660 then
	inst <= x"03DC0058";
end if;
if pc = 39664 then
	inst <= x"037E000C";
end if;
if pc = 39668 then
	inst <= x"C57DFFFC";
end if;
if pc = 39672 then
	inst <= x"82008034";
end if;
if pc = 39676 then
	inst <= x"07DC0058";
end if;
if pc = 39680 then
	inst <= x"82009B54";
end if;
if pc = 39684 then
	inst <= x"C04201DC";
end if;
if pc = 39688 then
	inst <= x"C8400014";
end if;
if pc = 39692 then
	inst <= x"C45C0050";
end if;
if pc = 39696 then
	inst <= x"CC3C0048";
end if;
if pc = 39700 then
	inst <= x"C17DFFFC";
end if;
if pc = 39704 then
	inst <= x"40204000";
end if;
if pc = 39708 then
	inst <= x"03DC005C";
end if;
if pc = 39712 then
	inst <= x"037E000C";
end if;
if pc = 39716 then
	inst <= x"C57DFFFC";
end if;
if pc = 39720 then
	inst <= x"82000844";
end if;
if pc = 39724 then
	inst <= x"07DC005C";
end if;
if pc = 39728 then
	inst <= x"C85C0048";
end if;
if pc = 39732 then
	inst <= x"48242000";
end if;
if pc = 39736 then
	inst <= x"C03C0050";
end if;
if pc = 39740 then
	inst <= x"C17DFFFC";
end if;
if pc = 39744 then
	inst <= x"03DC005C";
end if;
if pc = 39748 then
	inst <= x"037E000C";
end if;
if pc = 39752 then
	inst <= x"C57DFFFC";
end if;
if pc = 39756 then
	inst <= x"82008034";
end if;
if pc = 39760 then
	inst <= x"07DC005C";
end if;
if pc = 39764 then
	inst <= x"02800074";
end if;
if pc = 39768 then
	inst <= x"C03C003C";
end if;
if pc = 39772 then
	inst <= x"C05C0038";
end if;
if pc = 39776 then
	inst <= x"C07C0034";
end if;
if pc = 39780 then
	inst <= x"C17DFFFC";
end if;
if pc = 39784 then
	inst <= x"03DC005C";
end if;
if pc = 39788 then
	inst <= x"037E000C";
end if;
if pc = 39792 then
	inst <= x"C57DFFFC";
end if;
if pc = 39796 then
	inst <= x"82008280";
end if;
if pc = 39800 then
	inst <= x"07DC005C";
end if;
if pc = 39804 then
	inst <= x"C03C002C";
end if;
if pc = 39808 then
	inst <= x"C0420014";
end if;
if pc = 39812 then
	inst <= x"C0440000";
end if;
if pc = 39816 then
	inst <= x"C07C0030";
end if;
if pc = 39820 then
	inst <= x"C8260000";
end if;
if pc = 39824 then
	inst <= x"CC240000";
end if;
if pc = 39828 then
	inst <= x"C8260004";
end if;
if pc = 39832 then
	inst <= x"CC240004";
end if;
if pc = 39836 then
	inst <= x"C8260008";
end if;
if pc = 39840 then
	inst <= x"CC240008";
end if;
if pc = 39844 then
	inst <= x"82009BA8";
end if;
if pc = 39848 then
	inst <= x"02400001";
end if;
if pc = 39852 then
	inst <= x"C03C002C";
end if;
if pc = 39856 then
	inst <= x"C17DFFFC";
end if;
if pc = 39860 then
	inst <= x"03DC005C";
end if;
if pc = 39864 then
	inst <= x"037E000C";
end if;
if pc = 39868 then
	inst <= x"C57DFFFC";
end if;
if pc = 39872 then
	inst <= x"8200952C";
end if;
if pc = 39876 then
	inst <= x"07DC005C";
end if;
if pc = 39880 then
	inst <= x"82009BCC";
end if;
if pc = 39884 then
	inst <= x"C03C0024";
end if;
if pc = 39888 then
	inst <= x"06420001";
end if;
if pc = 39892 then
	inst <= x"C03C0018";
end if;
if pc = 39896 then
	inst <= x"02220001";
end if;
if pc = 39900 then
	inst <= x"02600005";
end if;
if pc = 39904 then
	inst <= x"86269BEC";
end if;
if pc = 39908 then
	inst <= x"06620005";
end if;
if pc = 39912 then
	inst <= x"82009BF0";
end if;
if pc = 39916 then
	inst <= x"00620000";
end if;
if pc = 39920 then
	inst <= x"C83C0010";
end if;
if pc = 39924 then
	inst <= x"C85C0008";
end if;
if pc = 39928 then
	inst <= x"C87C0000";
end if;
if pc = 39932 then
	inst <= x"C03C0020";
end if;
if pc = 39936 then
	inst <= x"82009870";
end if;
if pc = 39940 then
	inst <= x"C1FDFFFC";
end if;
if pc = 39944 then
	inst <= x"02800308";
end if;
if pc = 39948 then
	inst <= x"C8280000";
end if;
if pc = 39952 then
	inst <= x"02800300";
end if;
if pc = 39956 then
	inst <= x"C0880004";
end if;
if pc = 39960 then
	inst <= x"04448000";
end if;
if pc = 39964 then
	inst <= x"58440000";
end if;
if pc = 39968 then
	inst <= x"48224000";
end if;
if pc = 39972 then
	inst <= x"02400330";
end if;
if pc = 39976 then
	inst <= x"C8440000";
end if;
if pc = 39980 then
	inst <= x"48424000";
end if;
if pc = 39984 then
	inst <= x"0280033C";
end if;
if pc = 39988 then
	inst <= x"C8680000";
end if;
if pc = 39992 then
	inst <= x"40446000";
end if;
if pc = 39996 then
	inst <= x"C8640004";
end if;
if pc = 40000 then
	inst <= x"48626000";
end if;
if pc = 40004 then
	inst <= x"C8880004";
end if;
if pc = 40008 then
	inst <= x"40668000";
end if;
if pc = 40012 then
	inst <= x"C8840008";
end if;
if pc = 40016 then
	inst <= x"48228000";
end if;
if pc = 40020 then
	inst <= x"C8880008";
end if;
if pc = 40024 then
	inst <= x"40228000";
end if;
if pc = 40028 then
	inst <= x"024002F8";
end if;
if pc = 40032 then
	inst <= x"C0440000";
end if;
if pc = 40036 then
	inst <= x"06440001";
end if;
if pc = 40040 then
	inst <= x"41E06000";
end if;
if pc = 40044 then
	inst <= x"40602000";
end if;
if pc = 40048 then
	inst <= x"40204000";
end if;
if pc = 40052 then
	inst <= x"4041E000";
end if;
if pc = 40056 then
	inst <= x"82009870";
end if;
if pc = 40060 then
	inst <= x"02C002F8";
end if;
if pc = 40064 then
	inst <= x"C0EC0000";
end if;
if pc = 40068 then
	inst <= x"862E9C8C";
end if;
if pc = 40072 then
	inst <= x"C1FDFFFC";
end if;
if pc = 40076 then
	inst <= x"02E002EC";
end if;
if pc = 40080 then
	inst <= x"23020220";
end if;
if pc = 40084 then
	inst <= x"D1090000";
end if;
if pc = 40088 then
	inst <= x"C1100000";
end if;
if pc = 40092 then
	inst <= x"C8300000";
end if;
if pc = 40096 then
	inst <= x"CC2E0000";
end if;
if pc = 40100 then
	inst <= x"C8300004";
end if;
if pc = 40104 then
	inst <= x"CC2E0004";
end if;
if pc = 40108 then
	inst <= x"C8300008";
end if;
if pc = 40112 then
	inst <= x"CC2E0008";
end if;
if pc = 40116 then
	inst <= x"03040001";
end if;
if pc = 40120 then
	inst <= x"C12C0004";
end if;
if pc = 40124 then
	inst <= x"87129CC8";
end if;
if pc = 40128 then
	inst <= x"03000000";
end if;
if pc = 40132 then
	inst <= x"82009CF8";
end if;
if pc = 40136 then
	inst <= x"86049CD4";
end if;
if pc = 40140 then
	inst <= x"03000000";
end if;
if pc = 40144 then
	inst <= x"82009CF8";
end if;
if pc = 40148 then
	inst <= x"03020001";
end if;
if pc = 40152 then
	inst <= x"C12C0000";
end if;
if pc = 40156 then
	inst <= x"87129CE8";
end if;
if pc = 40160 then
	inst <= x"03000000";
end if;
if pc = 40164 then
	inst <= x"82009CF8";
end if;
if pc = 40168 then
	inst <= x"86029CF4";
end if;
if pc = 40172 then
	inst <= x"03000000";
end if;
if pc = 40176 then
	inst <= x"82009CF8";
end if;
if pc = 40180 then
	inst <= x"03000001";
end if;
if pc = 40184 then
	inst <= x"C4BC0000";
end if;
if pc = 40188 then
	inst <= x"C47C0004";
end if;
if pc = 40192 then
	inst <= x"C45C0008";
end if;
if pc = 40196 then
	inst <= x"C49C000C";
end if;
if pc = 40200 then
	inst <= x"C4DC0010";
end if;
if pc = 40204 then
	inst <= x"C43C0014";
end if;
if pc = 40208 then
	inst <= x"C4FC0018";
end if;
if pc = 40212 then
	inst <= x"83009E4C";
end if;
if pc = 40216 then
	inst <= x"03000000";
end if;
if pc = 40220 then
	inst <= x"23220220";
end if;
if pc = 40224 then
	inst <= x"D1292000";
end if;
if pc = 40228 then
	inst <= x"C1520008";
end if;
if pc = 40232 then
	inst <= x"C1540000";
end if;
if pc = 40236 then
	inst <= x"87409E48";
end if;
if pc = 40240 then
	inst <= x"C1520008";
end if;
if pc = 40244 then
	inst <= x"C1540000";
end if;
if pc = 40248 then
	inst <= x"22C20220";
end if;
if pc = 40252 then
	inst <= x"D0C6C000";
end if;
if pc = 40256 then
	inst <= x"C0CC0008";
end if;
if pc = 40260 then
	inst <= x"C0CC0000";
end if;
if pc = 40264 then
	inst <= x"82D49D54";
end if;
if pc = 40268 then
	inst <= x"02C00000";
end if;
if pc = 40272 then
	inst <= x"82009DB4";
end if;
if pc = 40276 then
	inst <= x"22C20220";
end if;
if pc = 40280 then
	inst <= x"D0CAC000";
end if;
if pc = 40284 then
	inst <= x"C0CC0008";
end if;
if pc = 40288 then
	inst <= x"C0CC0000";
end if;
if pc = 40292 then
	inst <= x"82D49D70";
end if;
if pc = 40296 then
	inst <= x"02C00000";
end if;
if pc = 40300 then
	inst <= x"82009DB4";
end if;
if pc = 40304 then
	inst <= x"06C20001";
end if;
if pc = 40308 then
	inst <= x"22CC0220";
end if;
if pc = 40312 then
	inst <= x"D0C8C000";
end if;
if pc = 40316 then
	inst <= x"C0CC0008";
end if;
if pc = 40320 then
	inst <= x"C0CC0000";
end if;
if pc = 40324 then
	inst <= x"82D49D90";
end if;
if pc = 40328 then
	inst <= x"02C00000";
end if;
if pc = 40332 then
	inst <= x"82009DB4";
end if;
if pc = 40336 then
	inst <= x"02C20001";
end if;
if pc = 40340 then
	inst <= x"22CC0220";
end if;
if pc = 40344 then
	inst <= x"D0C8C000";
end if;
if pc = 40348 then
	inst <= x"C0CC0008";
end if;
if pc = 40352 then
	inst <= x"C0CC0000";
end if;
if pc = 40356 then
	inst <= x"82D49DB0";
end if;
if pc = 40360 then
	inst <= x"02C00000";
end if;
if pc = 40364 then
	inst <= x"82009DB4";
end if;
if pc = 40368 then
	inst <= x"02C00001";
end if;
if pc = 40372 then
	inst <= x"82C09E24";
end if;
if pc = 40376 then
	inst <= x"C0D2000C";
end if;
if pc = 40380 then
	inst <= x"C0CC0000";
end if;
if pc = 40384 then
	inst <= x"82C09DF0";
end if;
if pc = 40388 then
	inst <= x"C17DFFFC";
end if;
if pc = 40392 then
	inst <= x"00460000";
end if;
if pc = 40396 then
	inst <= x"00680000";
end if;
if pc = 40400 then
	inst <= x"008A0000";
end if;
if pc = 40404 then
	inst <= x"00B00000";
end if;
if pc = 40408 then
	inst <= x"03DC0024";
end if;
if pc = 40412 then
	inst <= x"037E000C";
end if;
if pc = 40416 then
	inst <= x"C57DFFFC";
end if;
if pc = 40420 then
	inst <= x"82008F34";
end if;
if pc = 40424 then
	inst <= x"07DC0024";
end if;
if pc = 40428 then
	inst <= x"82009DF0";
end if;
if pc = 40432 then
	inst <= x"02C00001";
end if;
if pc = 40436 then
	inst <= x"C03C0014";
end if;
if pc = 40440 then
	inst <= x"C05C0008";
end if;
if pc = 40444 then
	inst <= x"C07C0004";
end if;
if pc = 40448 then
	inst <= x"C09C000C";
end if;
if pc = 40452 then
	inst <= x"C0BC0000";
end if;
if pc = 40456 then
	inst <= x"C17DFFFC";
end if;
if pc = 40460 then
	inst <= x"03DC0024";
end if;
if pc = 40464 then
	inst <= x"037E000C";
end if;
if pc = 40468 then
	inst <= x"C57DFFFC";
end if;
if pc = 40472 then
	inst <= x"8200925C";
end if;
if pc = 40476 then
	inst <= x"07DC0024";
end if;
if pc = 40480 then
	inst <= x"82009E44";
end if;
if pc = 40484 then
	inst <= x"C17DFFFC";
end if;
if pc = 40488 then
	inst <= x"00500000";
end if;
if pc = 40492 then
	inst <= x"00320000";
end if;
if pc = 40496 then
	inst <= x"03DC0024";
end if;
if pc = 40500 then
	inst <= x"037E000C";
end if;
if pc = 40504 then
	inst <= x"C57DFFFC";
end if;
if pc = 40508 then
	inst <= x"820090E0";
end if;
if pc = 40512 then
	inst <= x"07DC0024";
end if;
if pc = 40516 then
	inst <= x"82009E48";
end if;
if pc = 40520 then
	inst <= x"82009EBC";
end if;
if pc = 40524 then
	inst <= x"23020220";
end if;
if pc = 40528 then
	inst <= x"D1090000";
end if;
if pc = 40532 then
	inst <= x"03200000";
end if;
if pc = 40536 then
	inst <= x"C1500008";
end if;
if pc = 40540 then
	inst <= x"C1540000";
end if;
if pc = 40544 then
	inst <= x"87409EBC";
end if;
if pc = 40548 then
	inst <= x"C150000C";
end if;
if pc = 40552 then
	inst <= x"C1540000";
end if;
if pc = 40556 then
	inst <= x"C51C001C";
end if;
if pc = 40560 then
	inst <= x"83409E98";
end if;
if pc = 40564 then
	inst <= x"C17DFFFC";
end if;
if pc = 40568 then
	inst <= x"00520000";
end if;
if pc = 40572 then
	inst <= x"00300000";
end if;
if pc = 40576 then
	inst <= x"03DC0028";
end if;
if pc = 40580 then
	inst <= x"037E000C";
end if;
if pc = 40584 then
	inst <= x"C57DFFFC";
end if;
if pc = 40588 then
	inst <= x"8200874C";
end if;
if pc = 40592 then
	inst <= x"07DC0028";
end if;
if pc = 40596 then
	inst <= x"82009E98";
end if;
if pc = 40600 then
	inst <= x"02400001";
end if;
if pc = 40604 then
	inst <= x"C03C001C";
end if;
if pc = 40608 then
	inst <= x"C17DFFFC";
end if;
if pc = 40612 then
	inst <= x"03DC0028";
end if;
if pc = 40616 then
	inst <= x"037E000C";
end if;
if pc = 40620 then
	inst <= x"C57DFFFC";
end if;
if pc = 40624 then
	inst <= x"820090E0";
end if;
if pc = 40628 then
	inst <= x"07DC0028";
end if;
if pc = 40632 then
	inst <= x"82009EBC";
end if;
if pc = 40636 then
	inst <= x"C03C0018";
end if;
if pc = 40640 then
	inst <= x"C8220000";
end if;
if pc = 40644 then
	inst <= x"54420000";
end if;
if pc = 40648 then
	inst <= x"026000FF";
end if;
if pc = 40652 then
	inst <= x"86649EE0";
end if;
if pc = 40656 then
	inst <= x"86409ED8";
end if;
if pc = 40660 then
	inst <= x"82009EDC";
end if;
if pc = 40664 then
	inst <= x"02400000";
end if;
if pc = 40668 then
	inst <= x"82009EE4";
end if;
if pc = 40672 then
	inst <= x"024000FF";
end if;
if pc = 40676 then
	inst <= x"C17DFFFC";
end if;
if pc = 40680 then
	inst <= x"00240000";
end if;
if pc = 40684 then
	inst <= x"03DC0028";
end if;
if pc = 40688 then
	inst <= x"037E000C";
end if;
if pc = 40692 then
	inst <= x"C57DFFFC";
end if;
if pc = 40696 then
	inst <= x"8200078C";
end if;
if pc = 40700 then
	inst <= x"07DC0028";
end if;
if pc = 40704 then
	inst <= x"C03C0018";
end if;
if pc = 40708 then
	inst <= x"C8220004";
end if;
if pc = 40712 then
	inst <= x"54420000";
end if;
if pc = 40716 then
	inst <= x"026000FF";
end if;
if pc = 40720 then
	inst <= x"86649F24";
end if;
if pc = 40724 then
	inst <= x"86409F1C";
end if;
if pc = 40728 then
	inst <= x"82009F20";
end if;
if pc = 40732 then
	inst <= x"02400000";
end if;
if pc = 40736 then
	inst <= x"82009F28";
end if;
if pc = 40740 then
	inst <= x"024000FF";
end if;
if pc = 40744 then
	inst <= x"C17DFFFC";
end if;
if pc = 40748 then
	inst <= x"00240000";
end if;
if pc = 40752 then
	inst <= x"03DC0028";
end if;
if pc = 40756 then
	inst <= x"037E000C";
end if;
if pc = 40760 then
	inst <= x"C57DFFFC";
end if;
if pc = 40764 then
	inst <= x"8200078C";
end if;
if pc = 40768 then
	inst <= x"07DC0028";
end if;
if pc = 40772 then
	inst <= x"C03C0018";
end if;
if pc = 40776 then
	inst <= x"C8220008";
end if;
if pc = 40780 then
	inst <= x"54420000";
end if;
if pc = 40784 then
	inst <= x"026000FF";
end if;
if pc = 40788 then
	inst <= x"86649F68";
end if;
if pc = 40792 then
	inst <= x"86409F60";
end if;
if pc = 40796 then
	inst <= x"82009F64";
end if;
if pc = 40800 then
	inst <= x"02400000";
end if;
if pc = 40804 then
	inst <= x"82009F6C";
end if;
if pc = 40808 then
	inst <= x"024000FF";
end if;
if pc = 40812 then
	inst <= x"C17DFFFC";
end if;
if pc = 40816 then
	inst <= x"00240000";
end if;
if pc = 40820 then
	inst <= x"03DC0028";
end if;
if pc = 40824 then
	inst <= x"037E000C";
end if;
if pc = 40828 then
	inst <= x"C57DFFFC";
end if;
if pc = 40832 then
	inst <= x"8200078C";
end if;
if pc = 40836 then
	inst <= x"07DC0028";
end if;
if pc = 40840 then
	inst <= x"C03C0014";
end if;
if pc = 40844 then
	inst <= x"02220001";
end if;
if pc = 40848 then
	inst <= x"C05C0010";
end if;
if pc = 40852 then
	inst <= x"C0640000";
end if;
if pc = 40856 then
	inst <= x"86269FA0";
end if;
if pc = 40860 then
	inst <= x"C1FDFFFC";
end if;
if pc = 40864 then
	inst <= x"22620220";
end if;
if pc = 40868 then
	inst <= x"C09C000C";
end if;
if pc = 40872 then
	inst <= x"D0686000";
end if;
if pc = 40876 then
	inst <= x"C0660000";
end if;
if pc = 40880 then
	inst <= x"C8260000";
end if;
if pc = 40884 then
	inst <= x"C0BC0018";
end if;
if pc = 40888 then
	inst <= x"CC2A0000";
end if;
if pc = 40892 then
	inst <= x"C8260004";
end if;
if pc = 40896 then
	inst <= x"CC2A0004";
end if;
if pc = 40900 then
	inst <= x"C8260008";
end if;
if pc = 40904 then
	inst <= x"CC2A0008";
end if;
if pc = 40908 then
	inst <= x"C07C0008";
end if;
if pc = 40912 then
	inst <= x"02C60001";
end if;
if pc = 40916 then
	inst <= x"C0E40004";
end if;
if pc = 40920 then
	inst <= x"86CE9FE4";
end if;
if pc = 40924 then
	inst <= x"02400000";
end if;
if pc = 40928 then
	inst <= x"8200A014";
end if;
if pc = 40932 then
	inst <= x"86069FF0";
end if;
if pc = 40936 then
	inst <= x"02400000";
end if;
if pc = 40940 then
	inst <= x"8200A014";
end if;
if pc = 40944 then
	inst <= x"02C20001";
end if;
if pc = 40948 then
	inst <= x"C0440000";
end if;
if pc = 40952 then
	inst <= x"86C4A004";
end if;
if pc = 40956 then
	inst <= x"02400000";
end if;
if pc = 40960 then
	inst <= x"8200A014";
end if;
if pc = 40964 then
	inst <= x"8602A010";
end if;
if pc = 40968 then
	inst <= x"02400000";
end if;
if pc = 40972 then
	inst <= x"8200A014";
end if;
if pc = 40976 then
	inst <= x"02400001";
end if;
if pc = 40980 then
	inst <= x"C43C0020";
end if;
if pc = 40984 then
	inst <= x"8240A054";
end if;
if pc = 40988 then
	inst <= x"02C00000";
end if;
if pc = 40992 then
	inst <= x"C05C0004";
end if;
if pc = 40996 then
	inst <= x"C0FC0000";
end if;
if pc = 41000 then
	inst <= x"C17DFFFC";
end if;
if pc = 41004 then
	inst <= x"00AE0000";
end if;
if pc = 41008 then
	inst <= x"01260000";
end if;
if pc = 41012 then
	inst <= x"00640000";
end if;
if pc = 41016 then
	inst <= x"00520000";
end if;
if pc = 41020 then
	inst <= x"03DC002C";
end if;
if pc = 41024 then
	inst <= x"037E000C";
end if;
if pc = 41028 then
	inst <= x"C57DFFFC";
end if;
if pc = 41032 then
	inst <= x"8200925C";
end if;
if pc = 41036 then
	inst <= x"07DC002C";
end if;
if pc = 41040 then
	inst <= x"8200A080";
end if;
if pc = 41044 then
	inst <= x"22420220";
end if;
if pc = 41048 then
	inst <= x"D0484000";
end if;
if pc = 41052 then
	inst <= x"02C00000";
end if;
if pc = 41056 then
	inst <= x"C17DFFFC";
end if;
if pc = 41060 then
	inst <= x"00240000";
end if;
if pc = 41064 then
	inst <= x"004C0000";
end if;
if pc = 41068 then
	inst <= x"03DC002C";
end if;
if pc = 41072 then
	inst <= x"037E000C";
end if;
if pc = 41076 then
	inst <= x"C57DFFFC";
end if;
if pc = 41080 then
	inst <= x"820090E0";
end if;
if pc = 41084 then
	inst <= x"07DC002C";
end if;
if pc = 41088 then
	inst <= x"C03C0018";
end if;
if pc = 41092 then
	inst <= x"C8220000";
end if;
if pc = 41096 then
	inst <= x"54420000";
end if;
if pc = 41100 then
	inst <= x"026000FF";
end if;
if pc = 41104 then
	inst <= x"8664A0A4";
end if;
if pc = 41108 then
	inst <= x"8640A09C";
end if;
if pc = 41112 then
	inst <= x"8200A0A0";
end if;
if pc = 41116 then
	inst <= x"02400000";
end if;
if pc = 41120 then
	inst <= x"8200A0A8";
end if;
if pc = 41124 then
	inst <= x"024000FF";
end if;
if pc = 41128 then
	inst <= x"C17DFFFC";
end if;
if pc = 41132 then
	inst <= x"00240000";
end if;
if pc = 41136 then
	inst <= x"03DC002C";
end if;
if pc = 41140 then
	inst <= x"037E000C";
end if;
if pc = 41144 then
	inst <= x"C57DFFFC";
end if;
if pc = 41148 then
	inst <= x"8200078C";
end if;
if pc = 41152 then
	inst <= x"07DC002C";
end if;
if pc = 41156 then
	inst <= x"C03C0018";
end if;
if pc = 41160 then
	inst <= x"C8220004";
end if;
if pc = 41164 then
	inst <= x"54420000";
end if;
if pc = 41168 then
	inst <= x"026000FF";
end if;
if pc = 41172 then
	inst <= x"8664A0E8";
end if;
if pc = 41176 then
	inst <= x"8640A0E0";
end if;
if pc = 41180 then
	inst <= x"8200A0E4";
end if;
if pc = 41184 then
	inst <= x"02400000";
end if;
if pc = 41188 then
	inst <= x"8200A0EC";
end if;
if pc = 41192 then
	inst <= x"024000FF";
end if;
if pc = 41196 then
	inst <= x"C17DFFFC";
end if;
if pc = 41200 then
	inst <= x"00240000";
end if;
if pc = 41204 then
	inst <= x"03DC002C";
end if;
if pc = 41208 then
	inst <= x"037E000C";
end if;
if pc = 41212 then
	inst <= x"C57DFFFC";
end if;
if pc = 41216 then
	inst <= x"8200078C";
end if;
if pc = 41220 then
	inst <= x"07DC002C";
end if;
if pc = 41224 then
	inst <= x"C03C0018";
end if;
if pc = 41228 then
	inst <= x"C8220008";
end if;
if pc = 41232 then
	inst <= x"54220000";
end if;
if pc = 41236 then
	inst <= x"024000FF";
end if;
if pc = 41240 then
	inst <= x"8642A12C";
end if;
if pc = 41244 then
	inst <= x"8620A124";
end if;
if pc = 41248 then
	inst <= x"8200A128";
end if;
if pc = 41252 then
	inst <= x"02200000";
end if;
if pc = 41256 then
	inst <= x"8200A130";
end if;
if pc = 41260 then
	inst <= x"022000FF";
end if;
if pc = 41264 then
	inst <= x"C17DFFFC";
end if;
if pc = 41268 then
	inst <= x"03DC002C";
end if;
if pc = 41272 then
	inst <= x"037E000C";
end if;
if pc = 41276 then
	inst <= x"C57DFFFC";
end if;
if pc = 41280 then
	inst <= x"8200078C";
end if;
if pc = 41284 then
	inst <= x"07DC002C";
end if;
if pc = 41288 then
	inst <= x"C03C0020";
end if;
if pc = 41292 then
	inst <= x"02220001";
end if;
if pc = 41296 then
	inst <= x"C05C0008";
end if;
if pc = 41300 then
	inst <= x"C07C0004";
end if;
if pc = 41304 then
	inst <= x"C09C000C";
end if;
if pc = 41308 then
	inst <= x"C0BC0000";
end if;
if pc = 41312 then
	inst <= x"82009C7C";
end if;
if pc = 41316 then
	inst <= x"02C002F8";
end if;
if pc = 41320 then
	inst <= x"C0EC0004";
end if;
if pc = 41324 then
	inst <= x"862EA174";
end if;
if pc = 41328 then
	inst <= x"C1FDFFFC";
end if;
if pc = 41332 then
	inst <= x"C0EC0004";
end if;
if pc = 41336 then
	inst <= x"06EE0001";
end if;
if pc = 41340 then
	inst <= x"C4BC0000";
end if;
if pc = 41344 then
	inst <= x"C49C0004";
end if;
if pc = 41348 then
	inst <= x"C45C0008";
end if;
if pc = 41352 then
	inst <= x"C43C000C";
end if;
if pc = 41356 then
	inst <= x"C47C0010";
end if;
if pc = 41360 then
	inst <= x"C4DC0014";
end if;
if pc = 41364 then
	inst <= x"862EA19C";
end if;
if pc = 41368 then
	inst <= x"8200A1C4";
end if;
if pc = 41372 then
	inst <= x"02E20001";
end if;
if pc = 41376 then
	inst <= x"C17DFFFC";
end if;
if pc = 41380 then
	inst <= x"006A0000";
end if;
if pc = 41384 then
	inst <= x"004E0000";
end if;
if pc = 41388 then
	inst <= x"00280000";
end if;
if pc = 41392 then
	inst <= x"03DC0020";
end if;
if pc = 41396 then
	inst <= x"037E000C";
end if;
if pc = 41400 then
	inst <= x"C57DFFFC";
end if;
if pc = 41404 then
	inst <= x"82009C08";
end if;
if pc = 41408 then
	inst <= x"07DC0020";
end if;
if pc = 41412 then
	inst <= x"02200000";
end if;
if pc = 41416 then
	inst <= x"C05C0014";
end if;
if pc = 41420 then
	inst <= x"C0640000";
end if;
if pc = 41424 then
	inst <= x"8606A1D8";
end if;
if pc = 41428 then
	inst <= x"8200A390";
end if;
if pc = 41432 then
	inst <= x"026002EC";
end if;
if pc = 41436 then
	inst <= x"C09C0010";
end if;
if pc = 41440 then
	inst <= x"C0A80000";
end if;
if pc = 41444 then
	inst <= x"C0AA0000";
end if;
if pc = 41448 then
	inst <= x"C82A0000";
end if;
if pc = 41452 then
	inst <= x"CC260000";
end if;
if pc = 41456 then
	inst <= x"C82A0004";
end if;
if pc = 41460 then
	inst <= x"CC260004";
end if;
if pc = 41464 then
	inst <= x"C82A0008";
end if;
if pc = 41468 then
	inst <= x"CC260008";
end if;
if pc = 41472 then
	inst <= x"C0BC000C";
end if;
if pc = 41476 then
	inst <= x"02CA0001";
end if;
if pc = 41480 then
	inst <= x"C0E40004";
end if;
if pc = 41484 then
	inst <= x"86CEA218";
end if;
if pc = 41488 then
	inst <= x"02C00000";
end if;
if pc = 41492 then
	inst <= x"8200A23C";
end if;
if pc = 41496 then
	inst <= x"860AA224";
end if;
if pc = 41500 then
	inst <= x"02C00000";
end if;
if pc = 41504 then
	inst <= x"8200A23C";
end if;
if pc = 41508 then
	inst <= x"02C00001";
end if;
if pc = 41512 then
	inst <= x"C0E40000";
end if;
if pc = 41516 then
	inst <= x"86CEA238";
end if;
if pc = 41520 then
	inst <= x"02C00000";
end if;
if pc = 41524 then
	inst <= x"8200A23C";
end if;
if pc = 41528 then
	inst <= x"02C00001";
end if;
if pc = 41532 then
	inst <= x"C47C0018";
end if;
if pc = 41536 then
	inst <= x"82C0A278";
end if;
if pc = 41540 then
	inst <= x"02C00000";
end if;
if pc = 41544 then
	inst <= x"C0FC0008";
end if;
if pc = 41548 then
	inst <= x"C11C0004";
end if;
if pc = 41552 then
	inst <= x"C17DFFFC";
end if;
if pc = 41556 then
	inst <= x"006E0000";
end if;
if pc = 41560 then
	inst <= x"004A0000";
end if;
if pc = 41564 then
	inst <= x"00B00000";
end if;
if pc = 41568 then
	inst <= x"03DC0024";
end if;
if pc = 41572 then
	inst <= x"037E000C";
end if;
if pc = 41576 then
	inst <= x"C57DFFFC";
end if;
if pc = 41580 then
	inst <= x"8200925C";
end if;
if pc = 41584 then
	inst <= x"07DC0024";
end if;
if pc = 41588 then
	inst <= x"8200A29C";
end if;
if pc = 41592 then
	inst <= x"C0280000";
end if;
if pc = 41596 then
	inst <= x"02C00000";
end if;
if pc = 41600 then
	inst <= x"C17DFFFC";
end if;
if pc = 41604 then
	inst <= x"004C0000";
end if;
if pc = 41608 then
	inst <= x"03DC0024";
end if;
if pc = 41612 then
	inst <= x"037E000C";
end if;
if pc = 41616 then
	inst <= x"C57DFFFC";
end if;
if pc = 41620 then
	inst <= x"820090E0";
end if;
if pc = 41624 then
	inst <= x"07DC0024";
end if;
if pc = 41628 then
	inst <= x"C03C0018";
end if;
if pc = 41632 then
	inst <= x"C8220000";
end if;
if pc = 41636 then
	inst <= x"54420000";
end if;
if pc = 41640 then
	inst <= x"026000FF";
end if;
if pc = 41644 then
	inst <= x"8664A2C0";
end if;
if pc = 41648 then
	inst <= x"8640A2B8";
end if;
if pc = 41652 then
	inst <= x"8200A2BC";
end if;
if pc = 41656 then
	inst <= x"02400000";
end if;
if pc = 41660 then
	inst <= x"8200A2C4";
end if;
if pc = 41664 then
	inst <= x"024000FF";
end if;
if pc = 41668 then
	inst <= x"C17DFFFC";
end if;
if pc = 41672 then
	inst <= x"00240000";
end if;
if pc = 41676 then
	inst <= x"03DC0024";
end if;
if pc = 41680 then
	inst <= x"037E000C";
end if;
if pc = 41684 then
	inst <= x"C57DFFFC";
end if;
if pc = 41688 then
	inst <= x"8200078C";
end if;
if pc = 41692 then
	inst <= x"07DC0024";
end if;
if pc = 41696 then
	inst <= x"C03C0018";
end if;
if pc = 41700 then
	inst <= x"C8220004";
end if;
if pc = 41704 then
	inst <= x"54420000";
end if;
if pc = 41708 then
	inst <= x"026000FF";
end if;
if pc = 41712 then
	inst <= x"8664A304";
end if;
if pc = 41716 then
	inst <= x"8640A2FC";
end if;
if pc = 41720 then
	inst <= x"8200A300";
end if;
if pc = 41724 then
	inst <= x"02400000";
end if;
if pc = 41728 then
	inst <= x"8200A308";
end if;
if pc = 41732 then
	inst <= x"024000FF";
end if;
if pc = 41736 then
	inst <= x"C17DFFFC";
end if;
if pc = 41740 then
	inst <= x"00240000";
end if;
if pc = 41744 then
	inst <= x"03DC0024";
end if;
if pc = 41748 then
	inst <= x"037E000C";
end if;
if pc = 41752 then
	inst <= x"C57DFFFC";
end if;
if pc = 41756 then
	inst <= x"8200078C";
end if;
if pc = 41760 then
	inst <= x"07DC0024";
end if;
if pc = 41764 then
	inst <= x"C03C0018";
end if;
if pc = 41768 then
	inst <= x"C8220008";
end if;
if pc = 41772 then
	inst <= x"54220000";
end if;
if pc = 41776 then
	inst <= x"024000FF";
end if;
if pc = 41780 then
	inst <= x"8642A348";
end if;
if pc = 41784 then
	inst <= x"8620A340";
end if;
if pc = 41788 then
	inst <= x"8200A344";
end if;
if pc = 41792 then
	inst <= x"02200000";
end if;
if pc = 41796 then
	inst <= x"8200A34C";
end if;
if pc = 41800 then
	inst <= x"022000FF";
end if;
if pc = 41804 then
	inst <= x"C17DFFFC";
end if;
if pc = 41808 then
	inst <= x"03DC0024";
end if;
if pc = 41812 then
	inst <= x"037E000C";
end if;
if pc = 41816 then
	inst <= x"C57DFFFC";
end if;
if pc = 41820 then
	inst <= x"8200078C";
end if;
if pc = 41824 then
	inst <= x"07DC0024";
end if;
if pc = 41828 then
	inst <= x"02200001";
end if;
if pc = 41832 then
	inst <= x"C05C000C";
end if;
if pc = 41836 then
	inst <= x"C07C0008";
end if;
if pc = 41840 then
	inst <= x"C09C0010";
end if;
if pc = 41844 then
	inst <= x"C0BC0004";
end if;
if pc = 41848 then
	inst <= x"C17DFFFC";
end if;
if pc = 41852 then
	inst <= x"03DC0024";
end if;
if pc = 41856 then
	inst <= x"037E000C";
end if;
if pc = 41860 then
	inst <= x"C57DFFFC";
end if;
if pc = 41864 then
	inst <= x"82009C7C";
end if;
if pc = 41868 then
	inst <= x"07DC0024";
end if;
if pc = 41872 then
	inst <= x"C03C000C";
end if;
if pc = 41876 then
	inst <= x"02420001";
end if;
if pc = 41880 then
	inst <= x"C03C0000";
end if;
if pc = 41884 then
	inst <= x"02220002";
end if;
if pc = 41888 then
	inst <= x"02600005";
end if;
if pc = 41892 then
	inst <= x"8626A3B0";
end if;
if pc = 41896 then
	inst <= x"06620005";
end if;
if pc = 41900 then
	inst <= x"8200A3B4";
end if;
if pc = 41904 then
	inst <= x"00620000";
end if;
if pc = 41908 then
	inst <= x"C03C0014";
end if;
if pc = 41912 then
	inst <= x"C0820004";
end if;
if pc = 41916 then
	inst <= x"8648A3C4";
end if;
if pc = 41920 then
	inst <= x"8200A478";
end if;
if pc = 41924 then
	inst <= x"C0220004";
end if;
if pc = 41928 then
	inst <= x"06220001";
end if;
if pc = 41932 then
	inst <= x"C47C001C";
end if;
if pc = 41936 then
	inst <= x"C45C0020";
end if;
if pc = 41940 then
	inst <= x"8642A3DC";
end if;
if pc = 41944 then
	inst <= x"8200A404";
end if;
if pc = 41948 then
	inst <= x"02240001";
end if;
if pc = 41952 then
	inst <= x"C09C0008";
end if;
if pc = 41956 then
	inst <= x"C17DFFFC";
end if;
if pc = 41960 then
	inst <= x"00420000";
end if;
if pc = 41964 then
	inst <= x"00280000";
end if;
if pc = 41968 then
	inst <= x"03DC002C";
end if;
if pc = 41972 then
	inst <= x"037E000C";
end if;
if pc = 41976 then
	inst <= x"C57DFFFC";
end if;
if pc = 41980 then
	inst <= x"82009C08";
end if;
if pc = 41984 then
	inst <= x"07DC002C";
end if;
if pc = 41988 then
	inst <= x"02200000";
end if;
if pc = 41992 then
	inst <= x"C05C0020";
end if;
if pc = 41996 then
	inst <= x"C07C0010";
end if;
if pc = 42000 then
	inst <= x"C09C0004";
end if;
if pc = 42004 then
	inst <= x"C0BC0008";
end if;
if pc = 42008 then
	inst <= x"C17DFFFC";
end if;
if pc = 42012 then
	inst <= x"03DC002C";
end if;
if pc = 42016 then
	inst <= x"037E000C";
end if;
if pc = 42020 then
	inst <= x"C57DFFFC";
end if;
if pc = 42024 then
	inst <= x"82009C7C";
end if;
if pc = 42028 then
	inst <= x"07DC002C";
end if;
if pc = 42032 then
	inst <= x"C03C0020";
end if;
if pc = 42036 then
	inst <= x"02220001";
end if;
if pc = 42040 then
	inst <= x"C05C001C";
end if;
if pc = 42044 then
	inst <= x"02440002";
end if;
if pc = 42048 then
	inst <= x"02600005";
end if;
if pc = 42052 then
	inst <= x"8646A450";
end if;
if pc = 42056 then
	inst <= x"06A40005";
end if;
if pc = 42060 then
	inst <= x"8200A454";
end if;
if pc = 42064 then
	inst <= x"00A40000";
end if;
if pc = 42068 then
	inst <= x"C05C0004";
end if;
if pc = 42072 then
	inst <= x"C07C0008";
end if;
if pc = 42076 then
	inst <= x"C09C0010";
end if;
if pc = 42080 then
	inst <= x"C17DFFFC";
end if;
if pc = 42084 then
	inst <= x"03DC002C";
end if;
if pc = 42088 then
	inst <= x"037E000C";
end if;
if pc = 42092 then
	inst <= x"C57DFFFC";
end if;
if pc = 42096 then
	inst <= x"8200A164";
end if;
if pc = 42100 then
	inst <= x"07DC002C";
end if;
if pc = 42104 then
	inst <= x"C1FDFFFC";
end if;
if pc = 42108 then
	inst <= x"02200003";
end if;
if pc = 42112 then
	inst <= x"40200000";
end if;
if pc = 42116 then
	inst <= x"CC3C0000";
end if;
if pc = 42120 then
	inst <= x"C17DFFFC";
end if;
if pc = 42124 then
	inst <= x"03DC0010";
end if;
if pc = 42128 then
	inst <= x"037E000C";
end if;
if pc = 42132 then
	inst <= x"C57DFFFC";
end if;
if pc = 42136 then
	inst <= x"8200081C";
end if;
if pc = 42140 then
	inst <= x"07DC0010";
end if;
if pc = 42144 then
	inst <= x"02400003";
end if;
if pc = 42148 then
	inst <= x"C83C0000";
end if;
if pc = 42152 then
	inst <= x"C43C0008";
end if;
if pc = 42156 then
	inst <= x"C17DFFFC";
end if;
if pc = 42160 then
	inst <= x"00240000";
end if;
if pc = 42164 then
	inst <= x"03DC0014";
end if;
if pc = 42168 then
	inst <= x"037E000C";
end if;
if pc = 42172 then
	inst <= x"C57DFFFC";
end if;
if pc = 42176 then
	inst <= x"8200081C";
end if;
if pc = 42180 then
	inst <= x"07DC0014";
end if;
if pc = 42184 then
	inst <= x"00420000";
end if;
if pc = 42188 then
	inst <= x"02200005";
end if;
if pc = 42192 then
	inst <= x"C17DFFFC";
end if;
if pc = 42196 then
	inst <= x"03DC0014";
end if;
if pc = 42200 then
	inst <= x"037E000C";
end if;
if pc = 42204 then
	inst <= x"C57DFFFC";
end if;
if pc = 42208 then
	inst <= x"8200081C";
end if;
if pc = 42212 then
	inst <= x"07DC0014";
end if;
if pc = 42216 then
	inst <= x"02400003";
end if;
if pc = 42220 then
	inst <= x"C83C0000";
end if;
if pc = 42224 then
	inst <= x"C43C000C";
end if;
if pc = 42228 then
	inst <= x"C17DFFFC";
end if;
if pc = 42232 then
	inst <= x"00240000";
end if;
if pc = 42236 then
	inst <= x"03DC0018";
end if;
if pc = 42240 then
	inst <= x"037E000C";
end if;
if pc = 42244 then
	inst <= x"C57DFFFC";
end if;
if pc = 42248 then
	inst <= x"8200081C";
end if;
if pc = 42252 then
	inst <= x"07DC0018";
end if;
if pc = 42256 then
	inst <= x"C05C000C";
end if;
if pc = 42260 then
	inst <= x"C4240004";
end if;
if pc = 42264 then
	inst <= x"02200003";
end if;
if pc = 42268 then
	inst <= x"C83C0000";
end if;
if pc = 42272 then
	inst <= x"C17DFFFC";
end if;
if pc = 42276 then
	inst <= x"03DC0018";
end if;
if pc = 42280 then
	inst <= x"037E000C";
end if;
if pc = 42284 then
	inst <= x"C57DFFFC";
end if;
if pc = 42288 then
	inst <= x"8200081C";
end if;
if pc = 42292 then
	inst <= x"07DC0018";
end if;
if pc = 42296 then
	inst <= x"C05C000C";
end if;
if pc = 42300 then
	inst <= x"C4240008";
end if;
if pc = 42304 then
	inst <= x"02200003";
end if;
if pc = 42308 then
	inst <= x"C83C0000";
end if;
if pc = 42312 then
	inst <= x"C17DFFFC";
end if;
if pc = 42316 then
	inst <= x"03DC0018";
end if;
if pc = 42320 then
	inst <= x"037E000C";
end if;
if pc = 42324 then
	inst <= x"C57DFFFC";
end if;
if pc = 42328 then
	inst <= x"8200081C";
end if;
if pc = 42332 then
	inst <= x"07DC0018";
end if;
if pc = 42336 then
	inst <= x"C05C000C";
end if;
if pc = 42340 then
	inst <= x"C424000C";
end if;
if pc = 42344 then
	inst <= x"02200003";
end if;
if pc = 42348 then
	inst <= x"C83C0000";
end if;
if pc = 42352 then
	inst <= x"C17DFFFC";
end if;
if pc = 42356 then
	inst <= x"03DC0018";
end if;
if pc = 42360 then
	inst <= x"037E000C";
end if;
if pc = 42364 then
	inst <= x"C57DFFFC";
end if;
if pc = 42368 then
	inst <= x"8200081C";
end if;
if pc = 42372 then
	inst <= x"07DC0018";
end if;
if pc = 42376 then
	inst <= x"C05C000C";
end if;
if pc = 42380 then
	inst <= x"C4240010";
end if;
if pc = 42384 then
	inst <= x"02200005";
end if;
if pc = 42388 then
	inst <= x"02600000";
end if;
if pc = 42392 then
	inst <= x"C17DFFFC";
end if;
if pc = 42396 then
	inst <= x"00460000";
end if;
if pc = 42400 then
	inst <= x"03DC0018";
end if;
if pc = 42404 then
	inst <= x"037E000C";
end if;
if pc = 42408 then
	inst <= x"C57DFFFC";
end if;
if pc = 42412 then
	inst <= x"8200081C";
end if;
if pc = 42416 then
	inst <= x"07DC0018";
end if;
if pc = 42420 then
	inst <= x"02400005";
end if;
if pc = 42424 then
	inst <= x"02600000";
end if;
if pc = 42428 then
	inst <= x"C43C0010";
end if;
if pc = 42432 then
	inst <= x"C17DFFFC";
end if;
if pc = 42436 then
	inst <= x"00240000";
end if;
if pc = 42440 then
	inst <= x"00460000";
end if;
if pc = 42444 then
	inst <= x"03DC001C";
end if;
if pc = 42448 then
	inst <= x"037E000C";
end if;
if pc = 42452 then
	inst <= x"C57DFFFC";
end if;
if pc = 42456 then
	inst <= x"8200081C";
end if;
if pc = 42460 then
	inst <= x"07DC001C";
end if;
if pc = 42464 then
	inst <= x"02400003";
end if;
if pc = 42468 then
	inst <= x"C83C0000";
end if;
if pc = 42472 then
	inst <= x"C43C0014";
end if;
if pc = 42476 then
	inst <= x"C17DFFFC";
end if;
if pc = 42480 then
	inst <= x"00240000";
end if;
if pc = 42484 then
	inst <= x"03DC0020";
end if;
if pc = 42488 then
	inst <= x"037E000C";
end if;
if pc = 42492 then
	inst <= x"C57DFFFC";
end if;
if pc = 42496 then
	inst <= x"8200081C";
end if;
if pc = 42500 then
	inst <= x"07DC0020";
end if;
if pc = 42504 then
	inst <= x"00420000";
end if;
if pc = 42508 then
	inst <= x"02200005";
end if;
if pc = 42512 then
	inst <= x"C17DFFFC";
end if;
if pc = 42516 then
	inst <= x"03DC0020";
end if;
if pc = 42520 then
	inst <= x"037E000C";
end if;
if pc = 42524 then
	inst <= x"C57DFFFC";
end if;
if pc = 42528 then
	inst <= x"8200081C";
end if;
if pc = 42532 then
	inst <= x"07DC0020";
end if;
if pc = 42536 then
	inst <= x"02400003";
end if;
if pc = 42540 then
	inst <= x"C83C0000";
end if;
if pc = 42544 then
	inst <= x"C43C0018";
end if;
if pc = 42548 then
	inst <= x"C17DFFFC";
end if;
if pc = 42552 then
	inst <= x"00240000";
end if;
if pc = 42556 then
	inst <= x"03DC0024";
end if;
if pc = 42560 then
	inst <= x"037E000C";
end if;
if pc = 42564 then
	inst <= x"C57DFFFC";
end if;
if pc = 42568 then
	inst <= x"8200081C";
end if;
if pc = 42572 then
	inst <= x"07DC0024";
end if;
if pc = 42576 then
	inst <= x"C05C0018";
end if;
if pc = 42580 then
	inst <= x"C4240004";
end if;
if pc = 42584 then
	inst <= x"02200003";
end if;
if pc = 42588 then
	inst <= x"C83C0000";
end if;
if pc = 42592 then
	inst <= x"C17DFFFC";
end if;
if pc = 42596 then
	inst <= x"03DC0024";
end if;
if pc = 42600 then
	inst <= x"037E000C";
end if;
if pc = 42604 then
	inst <= x"C57DFFFC";
end if;
if pc = 42608 then
	inst <= x"8200081C";
end if;
if pc = 42612 then
	inst <= x"07DC0024";
end if;
if pc = 42616 then
	inst <= x"C05C0018";
end if;
if pc = 42620 then
	inst <= x"C4240008";
end if;
if pc = 42624 then
	inst <= x"02200003";
end if;
if pc = 42628 then
	inst <= x"C83C0000";
end if;
if pc = 42632 then
	inst <= x"C17DFFFC";
end if;
if pc = 42636 then
	inst <= x"03DC0024";
end if;
if pc = 42640 then
	inst <= x"037E000C";
end if;
if pc = 42644 then
	inst <= x"C57DFFFC";
end if;
if pc = 42648 then
	inst <= x"8200081C";
end if;
if pc = 42652 then
	inst <= x"07DC0024";
end if;
if pc = 42656 then
	inst <= x"C05C0018";
end if;
if pc = 42660 then
	inst <= x"C424000C";
end if;
if pc = 42664 then
	inst <= x"02200003";
end if;
if pc = 42668 then
	inst <= x"C83C0000";
end if;
if pc = 42672 then
	inst <= x"C17DFFFC";
end if;
if pc = 42676 then
	inst <= x"03DC0024";
end if;
if pc = 42680 then
	inst <= x"037E000C";
end if;
if pc = 42684 then
	inst <= x"C57DFFFC";
end if;
if pc = 42688 then
	inst <= x"8200081C";
end if;
if pc = 42692 then
	inst <= x"07DC0024";
end if;
if pc = 42696 then
	inst <= x"C05C0018";
end if;
if pc = 42700 then
	inst <= x"C4240010";
end if;
if pc = 42704 then
	inst <= x"02200003";
end if;
if pc = 42708 then
	inst <= x"C83C0000";
end if;
if pc = 42712 then
	inst <= x"C17DFFFC";
end if;
if pc = 42716 then
	inst <= x"03DC0024";
end if;
if pc = 42720 then
	inst <= x"037E000C";
end if;
if pc = 42724 then
	inst <= x"C57DFFFC";
end if;
if pc = 42728 then
	inst <= x"8200081C";
end if;
if pc = 42732 then
	inst <= x"07DC0024";
end if;
if pc = 42736 then
	inst <= x"00420000";
end if;
if pc = 42740 then
	inst <= x"02200005";
end if;
if pc = 42744 then
	inst <= x"C17DFFFC";
end if;
if pc = 42748 then
	inst <= x"03DC0024";
end if;
if pc = 42752 then
	inst <= x"037E000C";
end if;
if pc = 42756 then
	inst <= x"C57DFFFC";
end if;
if pc = 42760 then
	inst <= x"8200081C";
end if;
if pc = 42764 then
	inst <= x"07DC0024";
end if;
if pc = 42768 then
	inst <= x"02400003";
end if;
if pc = 42772 then
	inst <= x"C83C0000";
end if;
if pc = 42776 then
	inst <= x"C43C001C";
end if;
if pc = 42780 then
	inst <= x"C17DFFFC";
end if;
if pc = 42784 then
	inst <= x"00240000";
end if;
if pc = 42788 then
	inst <= x"03DC0028";
end if;
if pc = 42792 then
	inst <= x"037E000C";
end if;
if pc = 42796 then
	inst <= x"C57DFFFC";
end if;
if pc = 42800 then
	inst <= x"8200081C";
end if;
if pc = 42804 then
	inst <= x"07DC0028";
end if;
if pc = 42808 then
	inst <= x"C05C001C";
end if;
if pc = 42812 then
	inst <= x"C4240004";
end if;
if pc = 42816 then
	inst <= x"02200003";
end if;
if pc = 42820 then
	inst <= x"C83C0000";
end if;
if pc = 42824 then
	inst <= x"C17DFFFC";
end if;
if pc = 42828 then
	inst <= x"03DC0028";
end if;
if pc = 42832 then
	inst <= x"037E000C";
end if;
if pc = 42836 then
	inst <= x"C57DFFFC";
end if;
if pc = 42840 then
	inst <= x"8200081C";
end if;
if pc = 42844 then
	inst <= x"07DC0028";
end if;
if pc = 42848 then
	inst <= x"C05C001C";
end if;
if pc = 42852 then
	inst <= x"C4240008";
end if;
if pc = 42856 then
	inst <= x"02200003";
end if;
if pc = 42860 then
	inst <= x"C83C0000";
end if;
if pc = 42864 then
	inst <= x"C17DFFFC";
end if;
if pc = 42868 then
	inst <= x"03DC0028";
end if;
if pc = 42872 then
	inst <= x"037E000C";
end if;
if pc = 42876 then
	inst <= x"C57DFFFC";
end if;
if pc = 42880 then
	inst <= x"8200081C";
end if;
if pc = 42884 then
	inst <= x"07DC0028";
end if;
if pc = 42888 then
	inst <= x"C05C001C";
end if;
if pc = 42892 then
	inst <= x"C424000C";
end if;
if pc = 42896 then
	inst <= x"02200003";
end if;
if pc = 42900 then
	inst <= x"C83C0000";
end if;
if pc = 42904 then
	inst <= x"C17DFFFC";
end if;
if pc = 42908 then
	inst <= x"03DC0028";
end if;
if pc = 42912 then
	inst <= x"037E000C";
end if;
if pc = 42916 then
	inst <= x"C57DFFFC";
end if;
if pc = 42920 then
	inst <= x"8200081C";
end if;
if pc = 42924 then
	inst <= x"07DC0028";
end if;
if pc = 42928 then
	inst <= x"C05C001C";
end if;
if pc = 42932 then
	inst <= x"C4240010";
end if;
if pc = 42936 then
	inst <= x"02200001";
end if;
if pc = 42940 then
	inst <= x"02600000";
end if;
if pc = 42944 then
	inst <= x"C17DFFFC";
end if;
if pc = 42948 then
	inst <= x"00460000";
end if;
if pc = 42952 then
	inst <= x"03DC0028";
end if;
if pc = 42956 then
	inst <= x"037E000C";
end if;
if pc = 42960 then
	inst <= x"C57DFFFC";
end if;
if pc = 42964 then
	inst <= x"8200081C";
end if;
if pc = 42968 then
	inst <= x"07DC0028";
end if;
if pc = 42972 then
	inst <= x"02400003";
end if;
if pc = 42976 then
	inst <= x"C83C0000";
end if;
if pc = 42980 then
	inst <= x"C43C0020";
end if;
if pc = 42984 then
	inst <= x"C17DFFFC";
end if;
if pc = 42988 then
	inst <= x"00240000";
end if;
if pc = 42992 then
	inst <= x"03DC002C";
end if;
if pc = 42996 then
	inst <= x"037E000C";
end if;
if pc = 43000 then
	inst <= x"C57DFFFC";
end if;
if pc = 43004 then
	inst <= x"8200081C";
end if;
if pc = 43008 then
	inst <= x"07DC002C";
end if;
if pc = 43012 then
	inst <= x"00420000";
end if;
if pc = 43016 then
	inst <= x"02200005";
end if;
if pc = 43020 then
	inst <= x"C17DFFFC";
end if;
if pc = 43024 then
	inst <= x"03DC002C";
end if;
if pc = 43028 then
	inst <= x"037E000C";
end if;
if pc = 43032 then
	inst <= x"C57DFFFC";
end if;
if pc = 43036 then
	inst <= x"8200081C";
end if;
if pc = 43040 then
	inst <= x"07DC002C";
end if;
if pc = 43044 then
	inst <= x"02400003";
end if;
if pc = 43048 then
	inst <= x"C83C0000";
end if;
if pc = 43052 then
	inst <= x"C43C0024";
end if;
if pc = 43056 then
	inst <= x"C17DFFFC";
end if;
if pc = 43060 then
	inst <= x"00240000";
end if;
if pc = 43064 then
	inst <= x"03DC0030";
end if;
if pc = 43068 then
	inst <= x"037E000C";
end if;
if pc = 43072 then
	inst <= x"C57DFFFC";
end if;
if pc = 43076 then
	inst <= x"8200081C";
end if;
if pc = 43080 then
	inst <= x"07DC0030";
end if;
if pc = 43084 then
	inst <= x"C05C0024";
end if;
if pc = 43088 then
	inst <= x"C4240004";
end if;
if pc = 43092 then
	inst <= x"02200003";
end if;
if pc = 43096 then
	inst <= x"C83C0000";
end if;
if pc = 43100 then
	inst <= x"C17DFFFC";
end if;
if pc = 43104 then
	inst <= x"03DC0030";
end if;
if pc = 43108 then
	inst <= x"037E000C";
end if;
if pc = 43112 then
	inst <= x"C57DFFFC";
end if;
if pc = 43116 then
	inst <= x"8200081C";
end if;
if pc = 43120 then
	inst <= x"07DC0030";
end if;
if pc = 43124 then
	inst <= x"C05C0024";
end if;
if pc = 43128 then
	inst <= x"C4240008";
end if;
if pc = 43132 then
	inst <= x"02200003";
end if;
if pc = 43136 then
	inst <= x"C83C0000";
end if;
if pc = 43140 then
	inst <= x"C17DFFFC";
end if;
if pc = 43144 then
	inst <= x"03DC0030";
end if;
if pc = 43148 then
	inst <= x"037E000C";
end if;
if pc = 43152 then
	inst <= x"C57DFFFC";
end if;
if pc = 43156 then
	inst <= x"8200081C";
end if;
if pc = 43160 then
	inst <= x"07DC0030";
end if;
if pc = 43164 then
	inst <= x"C05C0024";
end if;
if pc = 43168 then
	inst <= x"C424000C";
end if;
if pc = 43172 then
	inst <= x"02200003";
end if;
if pc = 43176 then
	inst <= x"C83C0000";
end if;
if pc = 43180 then
	inst <= x"C17DFFFC";
end if;
if pc = 43184 then
	inst <= x"03DC0030";
end if;
if pc = 43188 then
	inst <= x"037E000C";
end if;
if pc = 43192 then
	inst <= x"C57DFFFC";
end if;
if pc = 43196 then
	inst <= x"8200081C";
end if;
if pc = 43200 then
	inst <= x"07DC0030";
end if;
if pc = 43204 then
	inst <= x"C05C0024";
end if;
if pc = 43208 then
	inst <= x"C4240010";
end if;
if pc = 43212 then
	inst <= x"003A0000";
end if;
if pc = 43216 then
	inst <= x"03BA0020";
end if;
if pc = 43220 then
	inst <= x"C442001C";
end if;
if pc = 43224 then
	inst <= x"C05C0020";
end if;
if pc = 43228 then
	inst <= x"C4420018";
end if;
if pc = 43232 then
	inst <= x"C05C001C";
end if;
if pc = 43236 then
	inst <= x"C4420014";
end if;
if pc = 43240 then
	inst <= x"C05C0018";
end if;
if pc = 43244 then
	inst <= x"C4420010";
end if;
if pc = 43248 then
	inst <= x"C05C0014";
end if;
if pc = 43252 then
	inst <= x"C442000C";
end if;
if pc = 43256 then
	inst <= x"C05C0010";
end if;
if pc = 43260 then
	inst <= x"C4420008";
end if;
if pc = 43264 then
	inst <= x"C05C000C";
end if;
if pc = 43268 then
	inst <= x"C4420004";
end if;
if pc = 43272 then
	inst <= x"C05C0008";
end if;
if pc = 43276 then
	inst <= x"C4420000";
end if;
if pc = 43280 then
	inst <= x"C1FDFFFC";
end if;
if pc = 43284 then
	inst <= x"8640AE10";
end if;
if pc = 43288 then
	inst <= x"02600003";
end if;
if pc = 43292 then
	inst <= x"40200000";
end if;
if pc = 43296 then
	inst <= x"C43C0000";
end if;
if pc = 43300 then
	inst <= x"C45C0004";
end if;
if pc = 43304 then
	inst <= x"CC3C0008";
end if;
if pc = 43308 then
	inst <= x"C17DFFFC";
end if;
if pc = 43312 then
	inst <= x"00260000";
end if;
if pc = 43316 then
	inst <= x"03DC0018";
end if;
if pc = 43320 then
	inst <= x"037E000C";
end if;
if pc = 43324 then
	inst <= x"C57DFFFC";
end if;
if pc = 43328 then
	inst <= x"8200081C";
end if;
if pc = 43332 then
	inst <= x"07DC0018";
end if;
if pc = 43336 then
	inst <= x"02400003";
end if;
if pc = 43340 then
	inst <= x"C83C0008";
end if;
if pc = 43344 then
	inst <= x"C43C0010";
end if;
if pc = 43348 then
	inst <= x"C17DFFFC";
end if;
if pc = 43352 then
	inst <= x"00240000";
end if;
if pc = 43356 then
	inst <= x"03DC001C";
end if;
if pc = 43360 then
	inst <= x"037E000C";
end if;
if pc = 43364 then
	inst <= x"C57DFFFC";
end if;
if pc = 43368 then
	inst <= x"8200081C";
end if;
if pc = 43372 then
	inst <= x"07DC001C";
end if;
if pc = 43376 then
	inst <= x"00420000";
end if;
if pc = 43380 then
	inst <= x"02200005";
end if;
if pc = 43384 then
	inst <= x"C17DFFFC";
end if;
if pc = 43388 then
	inst <= x"03DC001C";
end if;
if pc = 43392 then
	inst <= x"037E000C";
end if;
if pc = 43396 then
	inst <= x"C57DFFFC";
end if;
if pc = 43400 then
	inst <= x"8200081C";
end if;
if pc = 43404 then
	inst <= x"07DC001C";
end if;
if pc = 43408 then
	inst <= x"02400003";
end if;
if pc = 43412 then
	inst <= x"C83C0008";
end if;
if pc = 43416 then
	inst <= x"C43C0014";
end if;
if pc = 43420 then
	inst <= x"C17DFFFC";
end if;
if pc = 43424 then
	inst <= x"00240000";
end if;
if pc = 43428 then
	inst <= x"03DC0020";
end if;
if pc = 43432 then
	inst <= x"037E000C";
end if;
if pc = 43436 then
	inst <= x"C57DFFFC";
end if;
if pc = 43440 then
	inst <= x"8200081C";
end if;
if pc = 43444 then
	inst <= x"07DC0020";
end if;
if pc = 43448 then
	inst <= x"C05C0014";
end if;
if pc = 43452 then
	inst <= x"C4240004";
end if;
if pc = 43456 then
	inst <= x"02200003";
end if;
if pc = 43460 then
	inst <= x"C83C0008";
end if;
if pc = 43464 then
	inst <= x"C17DFFFC";
end if;
if pc = 43468 then
	inst <= x"03DC0020";
end if;
if pc = 43472 then
	inst <= x"037E000C";
end if;
if pc = 43476 then
	inst <= x"C57DFFFC";
end if;
if pc = 43480 then
	inst <= x"8200081C";
end if;
if pc = 43484 then
	inst <= x"07DC0020";
end if;
if pc = 43488 then
	inst <= x"C05C0014";
end if;
if pc = 43492 then
	inst <= x"C4240008";
end if;
if pc = 43496 then
	inst <= x"02200003";
end if;
if pc = 43500 then
	inst <= x"C83C0008";
end if;
if pc = 43504 then
	inst <= x"C17DFFFC";
end if;
if pc = 43508 then
	inst <= x"03DC0020";
end if;
if pc = 43512 then
	inst <= x"037E000C";
end if;
if pc = 43516 then
	inst <= x"C57DFFFC";
end if;
if pc = 43520 then
	inst <= x"8200081C";
end if;
if pc = 43524 then
	inst <= x"07DC0020";
end if;
if pc = 43528 then
	inst <= x"C05C0014";
end if;
if pc = 43532 then
	inst <= x"C424000C";
end if;
if pc = 43536 then
	inst <= x"02200003";
end if;
if pc = 43540 then
	inst <= x"C83C0008";
end if;
if pc = 43544 then
	inst <= x"C17DFFFC";
end if;
if pc = 43548 then
	inst <= x"03DC0020";
end if;
if pc = 43552 then
	inst <= x"037E000C";
end if;
if pc = 43556 then
	inst <= x"C57DFFFC";
end if;
if pc = 43560 then
	inst <= x"8200081C";
end if;
if pc = 43564 then
	inst <= x"07DC0020";
end if;
if pc = 43568 then
	inst <= x"C05C0014";
end if;
if pc = 43572 then
	inst <= x"C4240010";
end if;
if pc = 43576 then
	inst <= x"02200005";
end if;
if pc = 43580 then
	inst <= x"02600000";
end if;
if pc = 43584 then
	inst <= x"C17DFFFC";
end if;
if pc = 43588 then
	inst <= x"00460000";
end if;
if pc = 43592 then
	inst <= x"03DC0020";
end if;
if pc = 43596 then
	inst <= x"037E000C";
end if;
if pc = 43600 then
	inst <= x"C57DFFFC";
end if;
if pc = 43604 then
	inst <= x"8200081C";
end if;
if pc = 43608 then
	inst <= x"07DC0020";
end if;
if pc = 43612 then
	inst <= x"02400005";
end if;
if pc = 43616 then
	inst <= x"02600000";
end if;
if pc = 43620 then
	inst <= x"C43C0018";
end if;
if pc = 43624 then
	inst <= x"C17DFFFC";
end if;
if pc = 43628 then
	inst <= x"00240000";
end if;
if pc = 43632 then
	inst <= x"00460000";
end if;
if pc = 43636 then
	inst <= x"03DC0024";
end if;
if pc = 43640 then
	inst <= x"037E000C";
end if;
if pc = 43644 then
	inst <= x"C57DFFFC";
end if;
if pc = 43648 then
	inst <= x"8200081C";
end if;
if pc = 43652 then
	inst <= x"07DC0024";
end if;
if pc = 43656 then
	inst <= x"02400003";
end if;
if pc = 43660 then
	inst <= x"C83C0008";
end if;
if pc = 43664 then
	inst <= x"C43C001C";
end if;
if pc = 43668 then
	inst <= x"C17DFFFC";
end if;
if pc = 43672 then
	inst <= x"00240000";
end if;
if pc = 43676 then
	inst <= x"03DC0028";
end if;
if pc = 43680 then
	inst <= x"037E000C";
end if;
if pc = 43684 then
	inst <= x"C57DFFFC";
end if;
if pc = 43688 then
	inst <= x"8200081C";
end if;
if pc = 43692 then
	inst <= x"07DC0028";
end if;
if pc = 43696 then
	inst <= x"00420000";
end if;
if pc = 43700 then
	inst <= x"02200005";
end if;
if pc = 43704 then
	inst <= x"C17DFFFC";
end if;
if pc = 43708 then
	inst <= x"03DC0028";
end if;
if pc = 43712 then
	inst <= x"037E000C";
end if;
if pc = 43716 then
	inst <= x"C57DFFFC";
end if;
if pc = 43720 then
	inst <= x"8200081C";
end if;
if pc = 43724 then
	inst <= x"07DC0028";
end if;
if pc = 43728 then
	inst <= x"02400003";
end if;
if pc = 43732 then
	inst <= x"C83C0008";
end if;
if pc = 43736 then
	inst <= x"C43C0020";
end if;
if pc = 43740 then
	inst <= x"C17DFFFC";
end if;
if pc = 43744 then
	inst <= x"00240000";
end if;
if pc = 43748 then
	inst <= x"03DC002C";
end if;
if pc = 43752 then
	inst <= x"037E000C";
end if;
if pc = 43756 then
	inst <= x"C57DFFFC";
end if;
if pc = 43760 then
	inst <= x"8200081C";
end if;
if pc = 43764 then
	inst <= x"07DC002C";
end if;
if pc = 43768 then
	inst <= x"C05C0020";
end if;
if pc = 43772 then
	inst <= x"C4240004";
end if;
if pc = 43776 then
	inst <= x"02200003";
end if;
if pc = 43780 then
	inst <= x"C83C0008";
end if;
if pc = 43784 then
	inst <= x"C17DFFFC";
end if;
if pc = 43788 then
	inst <= x"03DC002C";
end if;
if pc = 43792 then
	inst <= x"037E000C";
end if;
if pc = 43796 then
	inst <= x"C57DFFFC";
end if;
if pc = 43800 then
	inst <= x"8200081C";
end if;
if pc = 43804 then
	inst <= x"07DC002C";
end if;
if pc = 43808 then
	inst <= x"C05C0020";
end if;
if pc = 43812 then
	inst <= x"C4240008";
end if;
if pc = 43816 then
	inst <= x"02200003";
end if;
if pc = 43820 then
	inst <= x"C83C0008";
end if;
if pc = 43824 then
	inst <= x"C17DFFFC";
end if;
if pc = 43828 then
	inst <= x"03DC002C";
end if;
if pc = 43832 then
	inst <= x"037E000C";
end if;
if pc = 43836 then
	inst <= x"C57DFFFC";
end if;
if pc = 43840 then
	inst <= x"8200081C";
end if;
if pc = 43844 then
	inst <= x"07DC002C";
end if;
if pc = 43848 then
	inst <= x"C05C0020";
end if;
if pc = 43852 then
	inst <= x"C424000C";
end if;
if pc = 43856 then
	inst <= x"02200003";
end if;
if pc = 43860 then
	inst <= x"C83C0008";
end if;
if pc = 43864 then
	inst <= x"C17DFFFC";
end if;
if pc = 43868 then
	inst <= x"03DC002C";
end if;
if pc = 43872 then
	inst <= x"037E000C";
end if;
if pc = 43876 then
	inst <= x"C57DFFFC";
end if;
if pc = 43880 then
	inst <= x"8200081C";
end if;
if pc = 43884 then
	inst <= x"07DC002C";
end if;
if pc = 43888 then
	inst <= x"C05C0020";
end if;
if pc = 43892 then
	inst <= x"C4240010";
end if;
if pc = 43896 then
	inst <= x"02200003";
end if;
if pc = 43900 then
	inst <= x"C83C0008";
end if;
if pc = 43904 then
	inst <= x"C17DFFFC";
end if;
if pc = 43908 then
	inst <= x"03DC002C";
end if;
if pc = 43912 then
	inst <= x"037E000C";
end if;
if pc = 43916 then
	inst <= x"C57DFFFC";
end if;
if pc = 43920 then
	inst <= x"8200081C";
end if;
if pc = 43924 then
	inst <= x"07DC002C";
end if;
if pc = 43928 then
	inst <= x"00420000";
end if;
if pc = 43932 then
	inst <= x"02200005";
end if;
if pc = 43936 then
	inst <= x"C17DFFFC";
end if;
if pc = 43940 then
	inst <= x"03DC002C";
end if;
if pc = 43944 then
	inst <= x"037E000C";
end if;
if pc = 43948 then
	inst <= x"C57DFFFC";
end if;
if pc = 43952 then
	inst <= x"8200081C";
end if;
if pc = 43956 then
	inst <= x"07DC002C";
end if;
if pc = 43960 then
	inst <= x"02400003";
end if;
if pc = 43964 then
	inst <= x"C83C0008";
end if;
if pc = 43968 then
	inst <= x"C43C0024";
end if;
if pc = 43972 then
	inst <= x"C17DFFFC";
end if;
if pc = 43976 then
	inst <= x"00240000";
end if;
if pc = 43980 then
	inst <= x"03DC0030";
end if;
if pc = 43984 then
	inst <= x"037E000C";
end if;
if pc = 43988 then
	inst <= x"C57DFFFC";
end if;
if pc = 43992 then
	inst <= x"8200081C";
end if;
if pc = 43996 then
	inst <= x"07DC0030";
end if;
if pc = 44000 then
	inst <= x"C05C0024";
end if;
if pc = 44004 then
	inst <= x"C4240004";
end if;
if pc = 44008 then
	inst <= x"02200003";
end if;
if pc = 44012 then
	inst <= x"C83C0008";
end if;
if pc = 44016 then
	inst <= x"C17DFFFC";
end if;
if pc = 44020 then
	inst <= x"03DC0030";
end if;
if pc = 44024 then
	inst <= x"037E000C";
end if;
if pc = 44028 then
	inst <= x"C57DFFFC";
end if;
if pc = 44032 then
	inst <= x"8200081C";
end if;
if pc = 44036 then
	inst <= x"07DC0030";
end if;
if pc = 44040 then
	inst <= x"C05C0024";
end if;
if pc = 44044 then
	inst <= x"C4240008";
end if;
if pc = 44048 then
	inst <= x"02200003";
end if;
if pc = 44052 then
	inst <= x"C83C0008";
end if;
if pc = 44056 then
	inst <= x"C17DFFFC";
end if;
if pc = 44060 then
	inst <= x"03DC0030";
end if;
if pc = 44064 then
	inst <= x"037E000C";
end if;
if pc = 44068 then
	inst <= x"C57DFFFC";
end if;
if pc = 44072 then
	inst <= x"8200081C";
end if;
if pc = 44076 then
	inst <= x"07DC0030";
end if;
if pc = 44080 then
	inst <= x"C05C0024";
end if;
if pc = 44084 then
	inst <= x"C424000C";
end if;
if pc = 44088 then
	inst <= x"02200003";
end if;
if pc = 44092 then
	inst <= x"C83C0008";
end if;
if pc = 44096 then
	inst <= x"C17DFFFC";
end if;
if pc = 44100 then
	inst <= x"03DC0030";
end if;
if pc = 44104 then
	inst <= x"037E000C";
end if;
if pc = 44108 then
	inst <= x"C57DFFFC";
end if;
if pc = 44112 then
	inst <= x"8200081C";
end if;
if pc = 44116 then
	inst <= x"07DC0030";
end if;
if pc = 44120 then
	inst <= x"C05C0024";
end if;
if pc = 44124 then
	inst <= x"C4240010";
end if;
if pc = 44128 then
	inst <= x"02200001";
end if;
if pc = 44132 then
	inst <= x"02600000";
end if;
if pc = 44136 then
	inst <= x"C17DFFFC";
end if;
if pc = 44140 then
	inst <= x"00460000";
end if;
if pc = 44144 then
	inst <= x"03DC0030";
end if;
if pc = 44148 then
	inst <= x"037E000C";
end if;
if pc = 44152 then
	inst <= x"C57DFFFC";
end if;
if pc = 44156 then
	inst <= x"8200081C";
end if;
if pc = 44160 then
	inst <= x"07DC0030";
end if;
if pc = 44164 then
	inst <= x"02400003";
end if;
if pc = 44168 then
	inst <= x"C83C0008";
end if;
if pc = 44172 then
	inst <= x"C43C0028";
end if;
if pc = 44176 then
	inst <= x"C17DFFFC";
end if;
if pc = 44180 then
	inst <= x"00240000";
end if;
if pc = 44184 then
	inst <= x"03DC0034";
end if;
if pc = 44188 then
	inst <= x"037E000C";
end if;
if pc = 44192 then
	inst <= x"C57DFFFC";
end if;
if pc = 44196 then
	inst <= x"8200081C";
end if;
if pc = 44200 then
	inst <= x"07DC0034";
end if;
if pc = 44204 then
	inst <= x"00420000";
end if;
if pc = 44208 then
	inst <= x"02200005";
end if;
if pc = 44212 then
	inst <= x"C17DFFFC";
end if;
if pc = 44216 then
	inst <= x"03DC0034";
end if;
if pc = 44220 then
	inst <= x"037E000C";
end if;
if pc = 44224 then
	inst <= x"C57DFFFC";
end if;
if pc = 44228 then
	inst <= x"8200081C";
end if;
if pc = 44232 then
	inst <= x"07DC0034";
end if;
if pc = 44236 then
	inst <= x"02400003";
end if;
if pc = 44240 then
	inst <= x"C83C0008";
end if;
if pc = 44244 then
	inst <= x"C43C002C";
end if;
if pc = 44248 then
	inst <= x"C17DFFFC";
end if;
if pc = 44252 then
	inst <= x"00240000";
end if;
if pc = 44256 then
	inst <= x"03DC0038";
end if;
if pc = 44260 then
	inst <= x"037E000C";
end if;
if pc = 44264 then
	inst <= x"C57DFFFC";
end if;
if pc = 44268 then
	inst <= x"8200081C";
end if;
if pc = 44272 then
	inst <= x"07DC0038";
end if;
if pc = 44276 then
	inst <= x"C05C002C";
end if;
if pc = 44280 then
	inst <= x"C4240004";
end if;
if pc = 44284 then
	inst <= x"02200003";
end if;
if pc = 44288 then
	inst <= x"C83C0008";
end if;
if pc = 44292 then
	inst <= x"C17DFFFC";
end if;
if pc = 44296 then
	inst <= x"03DC0038";
end if;
if pc = 44300 then
	inst <= x"037E000C";
end if;
if pc = 44304 then
	inst <= x"C57DFFFC";
end if;
if pc = 44308 then
	inst <= x"8200081C";
end if;
if pc = 44312 then
	inst <= x"07DC0038";
end if;
if pc = 44316 then
	inst <= x"C05C002C";
end if;
if pc = 44320 then
	inst <= x"C4240008";
end if;
if pc = 44324 then
	inst <= x"02200003";
end if;
if pc = 44328 then
	inst <= x"C83C0008";
end if;
if pc = 44332 then
	inst <= x"C17DFFFC";
end if;
if pc = 44336 then
	inst <= x"03DC0038";
end if;
if pc = 44340 then
	inst <= x"037E000C";
end if;
if pc = 44344 then
	inst <= x"C57DFFFC";
end if;
if pc = 44348 then
	inst <= x"8200081C";
end if;
if pc = 44352 then
	inst <= x"07DC0038";
end if;
if pc = 44356 then
	inst <= x"C05C002C";
end if;
if pc = 44360 then
	inst <= x"C424000C";
end if;
if pc = 44364 then
	inst <= x"02200003";
end if;
if pc = 44368 then
	inst <= x"C83C0008";
end if;
if pc = 44372 then
	inst <= x"C17DFFFC";
end if;
if pc = 44376 then
	inst <= x"03DC0038";
end if;
if pc = 44380 then
	inst <= x"037E000C";
end if;
if pc = 44384 then
	inst <= x"C57DFFFC";
end if;
if pc = 44388 then
	inst <= x"8200081C";
end if;
if pc = 44392 then
	inst <= x"07DC0038";
end if;
if pc = 44396 then
	inst <= x"C05C002C";
end if;
if pc = 44400 then
	inst <= x"C4240010";
end if;
if pc = 44404 then
	inst <= x"003A0000";
end if;
if pc = 44408 then
	inst <= x"03BA0020";
end if;
if pc = 44412 then
	inst <= x"C442001C";
end if;
if pc = 44416 then
	inst <= x"C05C0028";
end if;
if pc = 44420 then
	inst <= x"C4420018";
end if;
if pc = 44424 then
	inst <= x"C05C0024";
end if;
if pc = 44428 then
	inst <= x"C4420014";
end if;
if pc = 44432 then
	inst <= x"C05C0020";
end if;
if pc = 44436 then
	inst <= x"C4420010";
end if;
if pc = 44440 then
	inst <= x"C05C001C";
end if;
if pc = 44444 then
	inst <= x"C442000C";
end if;
if pc = 44448 then
	inst <= x"C05C0018";
end if;
if pc = 44452 then
	inst <= x"C4420008";
end if;
if pc = 44456 then
	inst <= x"C05C0014";
end if;
if pc = 44460 then
	inst <= x"C4420004";
end if;
if pc = 44464 then
	inst <= x"C05C0010";
end if;
if pc = 44468 then
	inst <= x"C4420000";
end if;
if pc = 44472 then
	inst <= x"C05C0004";
end if;
if pc = 44476 then
	inst <= x"22640220";
end if;
if pc = 44480 then
	inst <= x"C09C0000";
end if;
if pc = 44484 then
	inst <= x"D4286000";
end if;
if pc = 44488 then
	inst <= x"06240001";
end if;
if pc = 44492 then
	inst <= x"8620AE08";
end if;
if pc = 44496 then
	inst <= x"C43C0030";
end if;
if pc = 44500 then
	inst <= x"C17DFFFC";
end if;
if pc = 44504 then
	inst <= x"03DC003C";
end if;
if pc = 44508 then
	inst <= x"037E000C";
end if;
if pc = 44512 then
	inst <= x"C57DFFFC";
end if;
if pc = 44516 then
	inst <= x"8200A47C";
end if;
if pc = 44520 then
	inst <= x"07DC003C";
end if;
if pc = 44524 then
	inst <= x"C05C0030";
end if;
if pc = 44528 then
	inst <= x"22640220";
end if;
if pc = 44532 then
	inst <= x"C09C0000";
end if;
if pc = 44536 then
	inst <= x"D4286000";
end if;
if pc = 44540 then
	inst <= x"06440001";
end if;
if pc = 44544 then
	inst <= x"00280000";
end if;
if pc = 44548 then
	inst <= x"8200A914";
end if;
if pc = 44552 then
	inst <= x"00280000";
end if;
if pc = 44556 then
	inst <= x"C1FDFFFC";
end if;
if pc = 44560 then
	inst <= x"C1FDFFFC";
end if;
if pc = 44564 then
	inst <= x"02800005";
end if;
if pc = 44568 then
	inst <= x"8628AFA0";
end if;
if pc = 44572 then
	inst <= x"48622000";
end if;
if pc = 44576 then
	inst <= x"48844000";
end if;
if pc = 44580 then
	inst <= x"40668000";
end if;
if pc = 44584 then
	inst <= x"C88000A8";
end if;
if pc = 44588 then
	inst <= x"40668000";
end if;
if pc = 44592 then
	inst <= x"C47C0000";
end if;
if pc = 44596 then
	inst <= x"C45C0004";
end if;
if pc = 44600 then
	inst <= x"CC5C0008";
end if;
if pc = 44604 then
	inst <= x"CC3C0010";
end if;
if pc = 44608 then
	inst <= x"C17DFFFC";
end if;
if pc = 44612 then
	inst <= x"40206000";
end if;
if pc = 44616 then
	inst <= x"03DC0020";
end if;
if pc = 44620 then
	inst <= x"037E000C";
end if;
if pc = 44624 then
	inst <= x"C57DFFFC";
end if;
if pc = 44628 then
	inst <= x"8200083C";
end if;
if pc = 44632 then
	inst <= x"07DC0020";
end if;
if pc = 44636 then
	inst <= x"CC3C0018";
end if;
if pc = 44640 then
	inst <= x"C17DFFFC";
end if;
if pc = 44644 then
	inst <= x"03DC0028";
end if;
if pc = 44648 then
	inst <= x"037E000C";
end if;
if pc = 44652 then
	inst <= x"C57DFFFC";
end if;
if pc = 44656 then
	inst <= x"82000844";
end if;
if pc = 44660 then
	inst <= x"07DC0028";
end if;
if pc = 44664 then
	inst <= x"C85C0010";
end if;
if pc = 44668 then
	inst <= x"48242000";
end if;
if pc = 44672 then
	inst <= x"C85C0018";
end if;
if pc = 44676 then
	inst <= x"CC3C0020";
end if;
if pc = 44680 then
	inst <= x"C17DFFFC";
end if;
if pc = 44684 then
	inst <= x"40204000";
end if;
if pc = 44688 then
	inst <= x"03DC0030";
end if;
if pc = 44692 then
	inst <= x"037E000C";
end if;
if pc = 44696 then
	inst <= x"C57DFFFC";
end if;
if pc = 44700 then
	inst <= x"82000844";
end if;
if pc = 44704 then
	inst <= x"07DC0030";
end if;
if pc = 44708 then
	inst <= x"C85C0008";
end if;
if pc = 44712 then
	inst <= x"48242000";
end if;
if pc = 44716 then
	inst <= x"C85C0018";
end if;
if pc = 44720 then
	inst <= x"CC3C0028";
end if;
if pc = 44724 then
	inst <= x"C17DFFFC";
end if;
if pc = 44728 then
	inst <= x"40204000";
end if;
if pc = 44732 then
	inst <= x"03DC0038";
end if;
if pc = 44736 then
	inst <= x"037E000C";
end if;
if pc = 44740 then
	inst <= x"C57DFFFC";
end if;
if pc = 44744 then
	inst <= x"82000844";
end if;
if pc = 44748 then
	inst <= x"07DC0038";
end if;
if pc = 44752 then
	inst <= x"02200354";
end if;
if pc = 44756 then
	inst <= x"C05C0004";
end if;
if pc = 44760 then
	inst <= x"22440220";
end if;
if pc = 44764 then
	inst <= x"D0224000";
end if;
if pc = 44768 then
	inst <= x"C05C0000";
end if;
if pc = 44772 then
	inst <= x"22640220";
end if;
if pc = 44776 then
	inst <= x"D0626000";
end if;
if pc = 44780 then
	inst <= x"C0660000";
end if;
if pc = 44784 then
	inst <= x"C85C0020";
end if;
if pc = 44788 then
	inst <= x"CC460000";
end if;
if pc = 44792 then
	inst <= x"C87C0028";
end if;
if pc = 44796 then
	inst <= x"CC660004";
end if;
if pc = 44800 then
	inst <= x"CC260008";
end if;
if pc = 44804 then
	inst <= x"02640028";
end if;
if pc = 44808 then
	inst <= x"22660220";
end if;
if pc = 44812 then
	inst <= x"D0626000";
end if;
if pc = 44816 then
	inst <= x"C0660000";
end if;
if pc = 44820 then
	inst <= x"44806000";
end if;
if pc = 44824 then
	inst <= x"CC460000";
end if;
if pc = 44828 then
	inst <= x"CC260004";
end if;
if pc = 44832 then
	inst <= x"CC860008";
end if;
if pc = 44836 then
	inst <= x"02640050";
end if;
if pc = 44840 then
	inst <= x"22660220";
end if;
if pc = 44844 then
	inst <= x"D0626000";
end if;
if pc = 44848 then
	inst <= x"C0660000";
end if;
if pc = 44852 then
	inst <= x"44A04000";
end if;
if pc = 44856 then
	inst <= x"CC260000";
end if;
if pc = 44860 then
	inst <= x"CCA60004";
end if;
if pc = 44864 then
	inst <= x"CC860008";
end if;
if pc = 44868 then
	inst <= x"02640001";
end if;
if pc = 44872 then
	inst <= x"22660220";
end if;
if pc = 44876 then
	inst <= x"D0626000";
end if;
if pc = 44880 then
	inst <= x"C0660000";
end if;
if pc = 44884 then
	inst <= x"44202000";
end if;
if pc = 44888 then
	inst <= x"CCA60000";
end if;
if pc = 44892 then
	inst <= x"CC860004";
end if;
if pc = 44896 then
	inst <= x"CC260008";
end if;
if pc = 44900 then
	inst <= x"02640029";
end if;
if pc = 44904 then
	inst <= x"22660220";
end if;
if pc = 44908 then
	inst <= x"D0626000";
end if;
if pc = 44912 then
	inst <= x"C0660000";
end if;
if pc = 44916 then
	inst <= x"CCA60000";
end if;
if pc = 44920 then
	inst <= x"CC260004";
end if;
if pc = 44924 then
	inst <= x"CC660008";
end if;
if pc = 44928 then
	inst <= x"02440051";
end if;
if pc = 44932 then
	inst <= x"22440220";
end if;
if pc = 44936 then
	inst <= x"D0224000";
end if;
if pc = 44940 then
	inst <= x"C0220000";
end if;
if pc = 44944 then
	inst <= x"CC220000";
end if;
if pc = 44948 then
	inst <= x"CC420004";
end if;
if pc = 44952 then
	inst <= x"CC620008";
end if;
if pc = 44956 then
	inst <= x"C1FDFFFC";
end if;
if pc = 44960 then
	inst <= x"48244000";
end if;
if pc = 44964 then
	inst <= x"C840001C";
end if;
if pc = 44968 then
	inst <= x"40224000";
end if;
if pc = 44972 then
	inst <= x"C47C0000";
end if;
if pc = 44976 then
	inst <= x"C45C0004";
end if;
if pc = 44980 then
	inst <= x"CC9C0030";
end if;
if pc = 44984 then
	inst <= x"CC5C0038";
end if;
if pc = 44988 then
	inst <= x"C43C0040";
end if;
if pc = 44992 then
	inst <= x"CC7C0048";
end if;
if pc = 44996 then
	inst <= x"C17DFFFC";
end if;
if pc = 45000 then
	inst <= x"03DC0058";
end if;
if pc = 45004 then
	inst <= x"037E000C";
end if;
if pc = 45008 then
	inst <= x"C57DFFFC";
end if;
if pc = 45012 then
	inst <= x"8200083C";
end if;
if pc = 45016 then
	inst <= x"07DC0058";
end if;
if pc = 45020 then
	inst <= x"CC3C0050";
end if;
if pc = 45024 then
	inst <= x"C17DFFFC";
end if;
if pc = 45028 then
	inst <= x"03DC0060";
end if;
if pc = 45032 then
	inst <= x"037E000C";
end if;
if pc = 45036 then
	inst <= x"C57DFFFC";
end if;
if pc = 45040 then
	inst <= x"82000844";
end if;
if pc = 45044 then
	inst <= x"07DC0060";
end if;
if pc = 45048 then
	inst <= x"C8400068";
end if;
if pc = 45052 then
	inst <= x"48642000";
end if;
if pc = 45056 then
	inst <= x"C8800064";
end if;
if pc = 45060 then
	inst <= x"44668000";
end if;
if pc = 45064 then
	inst <= x"48662000";
end if;
if pc = 45068 then
	inst <= x"C8A00060";
end if;
if pc = 45072 then
	inst <= x"4466A000";
end if;
if pc = 45076 then
	inst <= x"48662000";
end if;
if pc = 45080 then
	inst <= x"C8C0005C";
end if;
if pc = 45084 then
	inst <= x"4066C000";
end if;
if pc = 45088 then
	inst <= x"48262000";
end if;
if pc = 45092 then
	inst <= x"C8600058";
end if;
if pc = 45096 then
	inst <= x"44226000";
end if;
if pc = 45100 then
	inst <= x"C8FC0048";
end if;
if pc = 45104 then
	inst <= x"4822E000";
end if;
if pc = 45108 then
	inst <= x"C9000098";
end if;
if pc = 45112 then
	inst <= x"CC7C0058";
end if;
if pc = 45116 then
	inst <= x"CCDC0060";
end if;
if pc = 45120 then
	inst <= x"CCBC0068";
end if;
if pc = 45124 then
	inst <= x"CC9C0070";
end if;
if pc = 45128 then
	inst <= x"CC5C0078";
end if;
if pc = 45132 then
	inst <= x"CD1C0080";
end if;
if pc = 45136 then
	inst <= x"CC3C0088";
end if;
if pc = 45140 then
	inst <= x"8E30B07C";
end if;
if pc = 45144 then
	inst <= x"45230000";
end if;
if pc = 45148 then
	inst <= x"C17DFFFC";
end if;
if pc = 45152 then
	inst <= x"40212000";
end if;
if pc = 45156 then
	inst <= x"03DC0098";
end if;
if pc = 45160 then
	inst <= x"037E000C";
end if;
if pc = 45164 then
	inst <= x"C57DFFFC";
end if;
if pc = 45168 then
	inst <= x"82000EC4";
end if;
if pc = 45172 then
	inst <= x"07DC0098";
end if;
if pc = 45176 then
	inst <= x"8200B0E8";
end if;
if pc = 45180 then
	inst <= x"8E02B0CC";
end if;
if pc = 45184 then
	inst <= x"C9200090";
end if;
if pc = 45188 then
	inst <= x"8F22B0AC";
end if;
if pc = 45192 then
	inst <= x"41230000";
end if;
if pc = 45196 then
	inst <= x"C17DFFFC";
end if;
if pc = 45200 then
	inst <= x"40212000";
end if;
if pc = 45204 then
	inst <= x"03DC0098";
end if;
if pc = 45208 then
	inst <= x"037E000C";
end if;
if pc = 45212 then
	inst <= x"C57DFFFC";
end if;
if pc = 45216 then
	inst <= x"82000EC4";
end if;
if pc = 45220 then
	inst <= x"07DC0098";
end if;
if pc = 45224 then
	inst <= x"8200B0C8";
end if;
if pc = 45228 then
	inst <= x"02200001";
end if;
if pc = 45232 then
	inst <= x"C17DFFFC";
end if;
if pc = 45236 then
	inst <= x"03DC0098";
end if;
if pc = 45240 then
	inst <= x"037E000C";
end if;
if pc = 45244 then
	inst <= x"C57DFFFC";
end if;
if pc = 45248 then
	inst <= x"8200084C";
end if;
if pc = 45252 then
	inst <= x"07DC0098";
end if;
if pc = 45256 then
	inst <= x"8200B0E8";
end if;
if pc = 45260 then
	inst <= x"0220FFFF";
end if;
if pc = 45264 then
	inst <= x"C17DFFFC";
end if;
if pc = 45268 then
	inst <= x"03DC0098";
end if;
if pc = 45272 then
	inst <= x"037E000C";
end if;
if pc = 45276 then
	inst <= x"C57DFFFC";
end if;
if pc = 45280 then
	inst <= x"8200084C";
end if;
if pc = 45284 then
	inst <= x"07DC0098";
end if;
if pc = 45288 then
	inst <= x"C85C0080";
end if;
if pc = 45292 then
	inst <= x"C87C0088";
end if;
if pc = 45296 then
	inst <= x"CC3C0090";
end if;
if pc = 45300 then
	inst <= x"8E64B11C";
end if;
if pc = 45304 then
	inst <= x"44664000";
end if;
if pc = 45308 then
	inst <= x"C17DFFFC";
end if;
if pc = 45312 then
	inst <= x"40206000";
end if;
if pc = 45316 then
	inst <= x"03DC00A0";
end if;
if pc = 45320 then
	inst <= x"037E000C";
end if;
if pc = 45324 then
	inst <= x"C57DFFFC";
end if;
if pc = 45328 then
	inst <= x"82001270";
end if;
if pc = 45332 then
	inst <= x"07DC00A0";
end if;
if pc = 45336 then
	inst <= x"8200B190";
end if;
if pc = 45340 then
	inst <= x"8E06B170";
end if;
if pc = 45344 then
	inst <= x"C8800090";
end if;
if pc = 45348 then
	inst <= x"8E86B14C";
end if;
if pc = 45352 then
	inst <= x"40664000";
end if;
if pc = 45356 then
	inst <= x"C17DFFFC";
end if;
if pc = 45360 then
	inst <= x"40206000";
end if;
if pc = 45364 then
	inst <= x"03DC00A0";
end if;
if pc = 45368 then
	inst <= x"037E000C";
end if;
if pc = 45372 then
	inst <= x"C57DFFFC";
end if;
if pc = 45376 then
	inst <= x"82001270";
end if;
if pc = 45380 then
	inst <= x"07DC00A0";
end if;
if pc = 45384 then
	inst <= x"8200B16C";
end if;
if pc = 45388 then
	inst <= x"02200001";
end if;
if pc = 45392 then
	inst <= x"C17DFFFC";
end if;
if pc = 45396 then
	inst <= x"40206000";
end if;
if pc = 45400 then
	inst <= x"03DC00A0";
end if;
if pc = 45404 then
	inst <= x"037E000C";
end if;
if pc = 45408 then
	inst <= x"C57DFFFC";
end if;
if pc = 45412 then
	inst <= x"82000B88";
end if;
if pc = 45416 then
	inst <= x"07DC00A0";
end if;
if pc = 45420 then
	inst <= x"8200B190";
end if;
if pc = 45424 then
	inst <= x"0220FFFF";
end if;
if pc = 45428 then
	inst <= x"C17DFFFC";
end if;
if pc = 45432 then
	inst <= x"40206000";
end if;
if pc = 45436 then
	inst <= x"03DC00A0";
end if;
if pc = 45440 then
	inst <= x"037E000C";
end if;
if pc = 45444 then
	inst <= x"C57DFFFC";
end if;
if pc = 45448 then
	inst <= x"82000B88";
end if;
if pc = 45452 then
	inst <= x"07DC00A0";
end if;
if pc = 45456 then
	inst <= x"C17DFFFC";
end if;
if pc = 45460 then
	inst <= x"03DC00A0";
end if;
if pc = 45464 then
	inst <= x"037E000C";
end if;
if pc = 45468 then
	inst <= x"C57DFFFC";
end if;
if pc = 45472 then
	inst <= x"82000844";
end if;
if pc = 45476 then
	inst <= x"07DC00A0";
end if;
if pc = 45480 then
	inst <= x"C85C0090";
end if;
if pc = 45484 then
	inst <= x"48242000";
end if;
if pc = 45488 then
	inst <= x"C85C0050";
end if;
if pc = 45492 then
	inst <= x"48224000";
end if;
if pc = 45496 then
	inst <= x"C03C0040";
end if;
if pc = 45500 then
	inst <= x"02220001";
end if;
if pc = 45504 then
	inst <= x"48422000";
end if;
if pc = 45508 then
	inst <= x"C87C0038";
end if;
if pc = 45512 then
	inst <= x"40446000";
end if;
if pc = 45516 then
	inst <= x"CC3C0098";
end if;
if pc = 45520 then
	inst <= x"C43C00A0";
end if;
if pc = 45524 then
	inst <= x"C17DFFFC";
end if;
if pc = 45528 then
	inst <= x"40204000";
end if;
if pc = 45532 then
	inst <= x"03DC00AC";
end if;
if pc = 45536 then
	inst <= x"037E000C";
end if;
if pc = 45540 then
	inst <= x"C57DFFFC";
end if;
if pc = 45544 then
	inst <= x"8200083C";
end if;
if pc = 45548 then
	inst <= x"07DC00AC";
end if;
if pc = 45552 then
	inst <= x"CC3C00A8";
end if;
if pc = 45556 then
	inst <= x"C17DFFFC";
end if;
if pc = 45560 then
	inst <= x"03DC00B8";
end if;
if pc = 45564 then
	inst <= x"037E000C";
end if;
if pc = 45568 then
	inst <= x"C57DFFFC";
end if;
if pc = 45572 then
	inst <= x"82000844";
end if;
if pc = 45576 then
	inst <= x"07DC00B8";
end if;
if pc = 45580 then
	inst <= x"C85C0078";
end if;
if pc = 45584 then
	inst <= x"48442000";
end if;
if pc = 45588 then
	inst <= x"C87C0070";
end if;
if pc = 45592 then
	inst <= x"44446000";
end if;
if pc = 45596 then
	inst <= x"48442000";
end if;
if pc = 45600 then
	inst <= x"C87C0068";
end if;
if pc = 45604 then
	inst <= x"44446000";
end if;
if pc = 45608 then
	inst <= x"48442000";
end if;
if pc = 45612 then
	inst <= x"C87C0060";
end if;
if pc = 45616 then
	inst <= x"40446000";
end if;
if pc = 45620 then
	inst <= x"48242000";
end if;
if pc = 45624 then
	inst <= x"C85C0058";
end if;
if pc = 45628 then
	inst <= x"44224000";
end if;
if pc = 45632 then
	inst <= x"C85C0030";
end if;
if pc = 45636 then
	inst <= x"48224000";
end if;
if pc = 45640 then
	inst <= x"C87C0080";
end if;
if pc = 45644 then
	inst <= x"CC3C00B0";
end if;
if pc = 45648 then
	inst <= x"8E26B278";
end if;
if pc = 45652 then
	inst <= x"44826000";
end if;
if pc = 45656 then
	inst <= x"C17DFFFC";
end if;
if pc = 45660 then
	inst <= x"40208000";
end if;
if pc = 45664 then
	inst <= x"03DC00C0";
end if;
if pc = 45668 then
	inst <= x"037E000C";
end if;
if pc = 45672 then
	inst <= x"C57DFFFC";
end if;
if pc = 45676 then
	inst <= x"82000EC4";
end if;
if pc = 45680 then
	inst <= x"07DC00C0";
end if;
if pc = 45684 then
	inst <= x"8200B2E4";
end if;
if pc = 45688 then
	inst <= x"8E02B2C8";
end if;
if pc = 45692 then
	inst <= x"C8800090";
end if;
if pc = 45696 then
	inst <= x"8E82B2A8";
end if;
if pc = 45700 then
	inst <= x"40826000";
end if;
if pc = 45704 then
	inst <= x"C17DFFFC";
end if;
if pc = 45708 then
	inst <= x"40208000";
end if;
if pc = 45712 then
	inst <= x"03DC00C0";
end if;
if pc = 45716 then
	inst <= x"037E000C";
end if;
if pc = 45720 then
	inst <= x"C57DFFFC";
end if;
if pc = 45724 then
	inst <= x"82000EC4";
end if;
if pc = 45728 then
	inst <= x"07DC00C0";
end if;
if pc = 45732 then
	inst <= x"8200B2C4";
end if;
if pc = 45736 then
	inst <= x"02200001";
end if;
if pc = 45740 then
	inst <= x"C17DFFFC";
end if;
if pc = 45744 then
	inst <= x"03DC00C0";
end if;
if pc = 45748 then
	inst <= x"037E000C";
end if;
if pc = 45752 then
	inst <= x"C57DFFFC";
end if;
if pc = 45756 then
	inst <= x"8200084C";
end if;
if pc = 45760 then
	inst <= x"07DC00C0";
end if;
if pc = 45764 then
	inst <= x"8200B2E4";
end if;
if pc = 45768 then
	inst <= x"0220FFFF";
end if;
if pc = 45772 then
	inst <= x"C17DFFFC";
end if;
if pc = 45776 then
	inst <= x"03DC00C0";
end if;
if pc = 45780 then
	inst <= x"037E000C";
end if;
if pc = 45784 then
	inst <= x"C57DFFFC";
end if;
if pc = 45788 then
	inst <= x"8200084C";
end if;
if pc = 45792 then
	inst <= x"07DC00C0";
end if;
if pc = 45796 then
	inst <= x"C85C0080";
end if;
if pc = 45800 then
	inst <= x"C87C00B0";
end if;
if pc = 45804 then
	inst <= x"CC3C00B8";
end if;
if pc = 45808 then
	inst <= x"8E64B318";
end if;
if pc = 45812 then
	inst <= x"44464000";
end if;
if pc = 45816 then
	inst <= x"C17DFFFC";
end if;
if pc = 45820 then
	inst <= x"40204000";
end if;
if pc = 45824 then
	inst <= x"03DC00C8";
end if;
if pc = 45828 then
	inst <= x"037E000C";
end if;
if pc = 45832 then
	inst <= x"C57DFFFC";
end if;
if pc = 45836 then
	inst <= x"82001270";
end if;
if pc = 45840 then
	inst <= x"07DC00C8";
end if;
if pc = 45844 then
	inst <= x"8200B38C";
end if;
if pc = 45848 then
	inst <= x"8E06B36C";
end if;
if pc = 45852 then
	inst <= x"C8800090";
end if;
if pc = 45856 then
	inst <= x"8E86B348";
end if;
if pc = 45860 then
	inst <= x"40464000";
end if;
if pc = 45864 then
	inst <= x"C17DFFFC";
end if;
if pc = 45868 then
	inst <= x"40204000";
end if;
if pc = 45872 then
	inst <= x"03DC00C8";
end if;
if pc = 45876 then
	inst <= x"037E000C";
end if;
if pc = 45880 then
	inst <= x"C57DFFFC";
end if;
if pc = 45884 then
	inst <= x"82001270";
end if;
if pc = 45888 then
	inst <= x"07DC00C8";
end if;
if pc = 45892 then
	inst <= x"8200B368";
end if;
if pc = 45896 then
	inst <= x"02200001";
end if;
if pc = 45900 then
	inst <= x"C17DFFFC";
end if;
if pc = 45904 then
	inst <= x"40206000";
end if;
if pc = 45908 then
	inst <= x"03DC00C8";
end if;
if pc = 45912 then
	inst <= x"037E000C";
end if;
if pc = 45916 then
	inst <= x"C57DFFFC";
end if;
if pc = 45920 then
	inst <= x"82000B88";
end if;
if pc = 45924 then
	inst <= x"07DC00C8";
end if;
if pc = 45928 then
	inst <= x"8200B38C";
end if;
if pc = 45932 then
	inst <= x"0220FFFF";
end if;
if pc = 45936 then
	inst <= x"C17DFFFC";
end if;
if pc = 45940 then
	inst <= x"40206000";
end if;
if pc = 45944 then
	inst <= x"03DC00C8";
end if;
if pc = 45948 then
	inst <= x"037E000C";
end if;
if pc = 45952 then
	inst <= x"C57DFFFC";
end if;
if pc = 45956 then
	inst <= x"82000B88";
end if;
if pc = 45960 then
	inst <= x"07DC00C8";
end if;
if pc = 45964 then
	inst <= x"C17DFFFC";
end if;
if pc = 45968 then
	inst <= x"03DC00C8";
end if;
if pc = 45972 then
	inst <= x"037E000C";
end if;
if pc = 45976 then
	inst <= x"C57DFFFC";
end if;
if pc = 45980 then
	inst <= x"82000844";
end if;
if pc = 45984 then
	inst <= x"07DC00C8";
end if;
if pc = 45988 then
	inst <= x"C85C00B8";
end if;
if pc = 45992 then
	inst <= x"48242000";
end if;
if pc = 45996 then
	inst <= x"C85C00A8";
end if;
if pc = 46000 then
	inst <= x"48424000";
end if;
if pc = 46004 then
	inst <= x"C83C0098";
end if;
if pc = 46008 then
	inst <= x"C87C0048";
end if;
if pc = 46012 then
	inst <= x"C89C0030";
end if;
if pc = 46016 then
	inst <= x"C03C00A0";
end if;
if pc = 46020 then
	inst <= x"C05C0004";
end if;
if pc = 46024 then
	inst <= x"C07C0000";
end if;
if pc = 46028 then
	inst <= x"8200AE14";
end if;
if pc = 46032 then
	inst <= x"8620B570";
end if;
if pc = 46036 then
	inst <= x"58420000";
end if;
if pc = 46040 then
	inst <= x"C8600010";
end if;
if pc = 46044 then
	inst <= x"48446000";
end if;
if pc = 46048 then
	inst <= x"C880000C";
end if;
if pc = 46052 then
	inst <= x"44A48000";
end if;
if pc = 46056 then
	inst <= x"02800000";
end if;
if pc = 46060 then
	inst <= x"40C00000";
end if;
if pc = 46064 then
	inst <= x"CC9C0000";
end if;
if pc = 46068 then
	inst <= x"CC7C0008";
end if;
if pc = 46072 then
	inst <= x"C43C0010";
end if;
if pc = 46076 then
	inst <= x"CC3C0018";
end if;
if pc = 46080 then
	inst <= x"CCDC0020";
end if;
if pc = 46084 then
	inst <= x"C45C0028";
end if;
if pc = 46088 then
	inst <= x"C47C002C";
end if;
if pc = 46092 then
	inst <= x"CC5C0030";
end if;
if pc = 46096 then
	inst <= x"C17DFFFC";
end if;
if pc = 46100 then
	inst <= x"00280000";
end if;
if pc = 46104 then
	inst <= x"40802000";
end if;
if pc = 46108 then
	inst <= x"4060A000";
end if;
if pc = 46112 then
	inst <= x"4040C000";
end if;
if pc = 46116 then
	inst <= x"4020C000";
end if;
if pc = 46120 then
	inst <= x"03DC0040";
end if;
if pc = 46124 then
	inst <= x"037E000C";
end if;
if pc = 46128 then
	inst <= x"C57DFFFC";
end if;
if pc = 46132 then
	inst <= x"8200AE14";
end if;
if pc = 46136 then
	inst <= x"07DC0040";
end if;
if pc = 46140 then
	inst <= x"C820001C";
end if;
if pc = 46144 then
	inst <= x"C85C0030";
end if;
if pc = 46148 then
	inst <= x"40642000";
end if;
if pc = 46152 then
	inst <= x"02200000";
end if;
if pc = 46156 then
	inst <= x"C05C002C";
end if;
if pc = 46160 then
	inst <= x"02640002";
end if;
if pc = 46164 then
	inst <= x"C85C0020";
end if;
if pc = 46168 then
	inst <= x"C89C0018";
end if;
if pc = 46172 then
	inst <= x"C09C0028";
end if;
if pc = 46176 then
	inst <= x"CC3C0038";
end if;
if pc = 46180 then
	inst <= x"C17DFFFC";
end if;
if pc = 46184 then
	inst <= x"00480000";
end if;
if pc = 46188 then
	inst <= x"40204000";
end if;
if pc = 46192 then
	inst <= x"03DC0048";
end if;
if pc = 46196 then
	inst <= x"037E000C";
end if;
if pc = 46200 then
	inst <= x"C57DFFFC";
end if;
if pc = 46204 then
	inst <= x"8200AE14";
end if;
if pc = 46208 then
	inst <= x"07DC0048";
end if;
if pc = 46212 then
	inst <= x"C03C0010";
end if;
if pc = 46216 then
	inst <= x"06220001";
end if;
if pc = 46220 then
	inst <= x"C05C0028";
end if;
if pc = 46224 then
	inst <= x"02440001";
end if;
if pc = 46228 then
	inst <= x"02600005";
end if;
if pc = 46232 then
	inst <= x"8646B4A4";
end if;
if pc = 46236 then
	inst <= x"06440005";
end if;
if pc = 46240 then
	inst <= x"8200B4A4";
end if;
if pc = 46244 then
	inst <= x"8620B56C";
end if;
if pc = 46248 then
	inst <= x"58220000";
end if;
if pc = 46252 then
	inst <= x"C85C0008";
end if;
if pc = 46256 then
	inst <= x"48224000";
end if;
if pc = 46260 then
	inst <= x"C85C0000";
end if;
if pc = 46264 then
	inst <= x"44624000";
end if;
if pc = 46268 then
	inst <= x"02600000";
end if;
if pc = 46272 then
	inst <= x"C85C0020";
end if;
if pc = 46276 then
	inst <= x"C89C0018";
end if;
if pc = 46280 then
	inst <= x"C09C002C";
end if;
if pc = 46284 then
	inst <= x"C43C0040";
end if;
if pc = 46288 then
	inst <= x"C45C0044";
end if;
if pc = 46292 then
	inst <= x"CC3C0048";
end if;
if pc = 46296 then
	inst <= x"C17DFFFC";
end if;
if pc = 46300 then
	inst <= x"00260000";
end if;
if pc = 46304 then
	inst <= x"00680000";
end if;
if pc = 46308 then
	inst <= x"40204000";
end if;
if pc = 46312 then
	inst <= x"03DC0058";
end if;
if pc = 46316 then
	inst <= x"037E000C";
end if;
if pc = 46320 then
	inst <= x"C57DFFFC";
end if;
if pc = 46324 then
	inst <= x"8200AE14";
end if;
if pc = 46328 then
	inst <= x"07DC0058";
end if;
if pc = 46332 then
	inst <= x"C83C0038";
end if;
if pc = 46336 then
	inst <= x"C85C0048";
end if;
if pc = 46340 then
	inst <= x"40642000";
end if;
if pc = 46344 then
	inst <= x"02200000";
end if;
if pc = 46348 then
	inst <= x"C05C002C";
end if;
if pc = 46352 then
	inst <= x"02640002";
end if;
if pc = 46356 then
	inst <= x"C83C0020";
end if;
if pc = 46360 then
	inst <= x"C89C0018";
end if;
if pc = 46364 then
	inst <= x"C09C0044";
end if;
if pc = 46368 then
	inst <= x"C17DFFFC";
end if;
if pc = 46372 then
	inst <= x"00480000";
end if;
if pc = 46376 then
	inst <= x"40402000";
end if;
if pc = 46380 then
	inst <= x"03DC0058";
end if;
if pc = 46384 then
	inst <= x"037E000C";
end if;
if pc = 46388 then
	inst <= x"C57DFFFC";
end if;
if pc = 46392 then
	inst <= x"8200AE14";
end if;
if pc = 46396 then
	inst <= x"07DC0058";
end if;
if pc = 46400 then
	inst <= x"C03C0040";
end if;
if pc = 46404 then
	inst <= x"06220001";
end if;
if pc = 46408 then
	inst <= x"C05C0044";
end if;
if pc = 46412 then
	inst <= x"02440001";
end if;
if pc = 46416 then
	inst <= x"02600005";
end if;
if pc = 46420 then
	inst <= x"8646B560";
end if;
if pc = 46424 then
	inst <= x"06440005";
end if;
if pc = 46428 then
	inst <= x"8200B560";
end if;
if pc = 46432 then
	inst <= x"C83C0018";
end if;
if pc = 46436 then
	inst <= x"C07C002C";
end if;
if pc = 46440 then
	inst <= x"8200B3D0";
end if;
if pc = 46444 then
	inst <= x"C1FDFFFC";
end if;
if pc = 46448 then
	inst <= x"C1FDFFFC";
end if;
if pc = 46452 then
	inst <= x"8620B6F8";
end if;
if pc = 46456 then
	inst <= x"58220000";
end if;
if pc = 46460 then
	inst <= x"C8400010";
end if;
if pc = 46464 then
	inst <= x"48224000";
end if;
if pc = 46468 then
	inst <= x"C860000C";
end if;
if pc = 46472 then
	inst <= x"44826000";
end if;
if pc = 46476 then
	inst <= x"C8200008";
end if;
if pc = 46480 then
	inst <= x"02800000";
end if;
if pc = 46484 then
	inst <= x"40A00000";
end if;
if pc = 46488 then
	inst <= x"CC5C0000";
end if;
if pc = 46492 then
	inst <= x"C43C0008";
end if;
if pc = 46496 then
	inst <= x"CC9C0010";
end if;
if pc = 46500 then
	inst <= x"CC7C0018";
end if;
if pc = 46504 then
	inst <= x"CCBC0020";
end if;
if pc = 46508 then
	inst <= x"C45C0028";
end if;
if pc = 46512 then
	inst <= x"C47C002C";
end if;
if pc = 46516 then
	inst <= x"C17DFFFC";
end if;
if pc = 46520 then
	inst <= x"00280000";
end if;
if pc = 46524 then
	inst <= x"40602000";
end if;
if pc = 46528 then
	inst <= x"4040A000";
end if;
if pc = 46532 then
	inst <= x"4020A000";
end if;
if pc = 46536 then
	inst <= x"03DC0038";
end if;
if pc = 46540 then
	inst <= x"037E000C";
end if;
if pc = 46544 then
	inst <= x"C57DFFFC";
end if;
if pc = 46548 then
	inst <= x"8200AE14";
end if;
if pc = 46552 then
	inst <= x"07DC0038";
end if;
if pc = 46556 then
	inst <= x"02200000";
end if;
if pc = 46560 then
	inst <= x"C05C002C";
end if;
if pc = 46564 then
	inst <= x"02640002";
end if;
if pc = 46568 then
	inst <= x"C83C0020";
end if;
if pc = 46572 then
	inst <= x"C87C0018";
end if;
if pc = 46576 then
	inst <= x"C89C0010";
end if;
if pc = 46580 then
	inst <= x"C09C0028";
end if;
if pc = 46584 then
	inst <= x"C17DFFFC";
end if;
if pc = 46588 then
	inst <= x"00480000";
end if;
if pc = 46592 then
	inst <= x"40402000";
end if;
if pc = 46596 then
	inst <= x"03DC0038";
end if;
if pc = 46600 then
	inst <= x"037E000C";
end if;
if pc = 46604 then
	inst <= x"C57DFFFC";
end if;
if pc = 46608 then
	inst <= x"8200AE14";
end if;
if pc = 46612 then
	inst <= x"07DC0038";
end if;
if pc = 46616 then
	inst <= x"02200003";
end if;
if pc = 46620 then
	inst <= x"C05C0028";
end if;
if pc = 46624 then
	inst <= x"02640001";
end if;
if pc = 46628 then
	inst <= x"02800005";
end if;
if pc = 46632 then
	inst <= x"8668B634";
end if;
if pc = 46636 then
	inst <= x"06660005";
end if;
if pc = 46640 then
	inst <= x"8200B634";
end if;
if pc = 46644 then
	inst <= x"C83C0010";
end if;
if pc = 46648 then
	inst <= x"C09C002C";
end if;
if pc = 46652 then
	inst <= x"C17DFFFC";
end if;
if pc = 46656 then
	inst <= x"00460000";
end if;
if pc = 46660 then
	inst <= x"00680000";
end if;
if pc = 46664 then
	inst <= x"03DC0038";
end if;
if pc = 46668 then
	inst <= x"037E000C";
end if;
if pc = 46672 then
	inst <= x"C57DFFFC";
end if;
if pc = 46676 then
	inst <= x"8200B3D0";
end if;
if pc = 46680 then
	inst <= x"07DC0038";
end if;
if pc = 46684 then
	inst <= x"C03C0008";
end if;
if pc = 46688 then
	inst <= x"06220001";
end if;
if pc = 46692 then
	inst <= x"C05C0028";
end if;
if pc = 46696 then
	inst <= x"02440002";
end if;
if pc = 46700 then
	inst <= x"02600005";
end if;
if pc = 46704 then
	inst <= x"8646B67C";
end if;
if pc = 46708 then
	inst <= x"06440005";
end if;
if pc = 46712 then
	inst <= x"8200B67C";
end if;
if pc = 46716 then
	inst <= x"C07C002C";
end if;
if pc = 46720 then
	inst <= x"02660004";
end if;
if pc = 46724 then
	inst <= x"8620B6F4";
end if;
if pc = 46728 then
	inst <= x"58220000";
end if;
if pc = 46732 then
	inst <= x"C85C0000";
end if;
if pc = 46736 then
	inst <= x"48224000";
end if;
if pc = 46740 then
	inst <= x"C85C0018";
end if;
if pc = 46744 then
	inst <= x"44224000";
end if;
if pc = 46748 then
	inst <= x"02800004";
end if;
if pc = 46752 then
	inst <= x"C47C0030";
end if;
if pc = 46756 then
	inst <= x"C45C0034";
end if;
if pc = 46760 then
	inst <= x"C43C0038";
end if;
if pc = 46764 then
	inst <= x"C17DFFFC";
end if;
if pc = 46768 then
	inst <= x"00280000";
end if;
if pc = 46772 then
	inst <= x"03DC0044";
end if;
if pc = 46776 then
	inst <= x"037E000C";
end if;
if pc = 46780 then
	inst <= x"C57DFFFC";
end if;
if pc = 46784 then
	inst <= x"8200B3D0";
end if;
if pc = 46788 then
	inst <= x"07DC0044";
end if;
if pc = 46792 then
	inst <= x"C03C0038";
end if;
if pc = 46796 then
	inst <= x"06220001";
end if;
if pc = 46800 then
	inst <= x"C05C0034";
end if;
if pc = 46804 then
	inst <= x"02440002";
end if;
if pc = 46808 then
	inst <= x"02600005";
end if;
if pc = 46812 then
	inst <= x"8646B6E8";
end if;
if pc = 46816 then
	inst <= x"06440005";
end if;
if pc = 46820 then
	inst <= x"8200B6E8";
end if;
if pc = 46824 then
	inst <= x"C07C0030";
end if;
if pc = 46828 then
	inst <= x"02660004";
end if;
if pc = 46832 then
	inst <= x"8200B574";
end if;
if pc = 46836 then
	inst <= x"C1FDFFFC";
end if;
if pc = 46840 then
	inst <= x"C1FDFFFC";
end if;
if pc = 46844 then
	inst <= x"8640B928";
end if;
if pc = 46848 then
	inst <= x"02600003";
end if;
if pc = 46852 then
	inst <= x"40200000";
end if;
if pc = 46856 then
	inst <= x"CC3C0000";
end if;
if pc = 46860 then
	inst <= x"C43C0008";
end if;
if pc = 46864 then
	inst <= x"C45C000C";
end if;
if pc = 46868 then
	inst <= x"C17DFFFC";
end if;
if pc = 46872 then
	inst <= x"00260000";
end if;
if pc = 46876 then
	inst <= x"03DC0018";
end if;
if pc = 46880 then
	inst <= x"037E000C";
end if;
if pc = 46884 then
	inst <= x"C57DFFFC";
end if;
if pc = 46888 then
	inst <= x"8200081C";
end if;
if pc = 46892 then
	inst <= x"07DC0018";
end if;
if pc = 46896 then
	inst <= x"00420000";
end if;
if pc = 46900 then
	inst <= x"022000C4";
end if;
if pc = 46904 then
	inst <= x"C0620000";
end if;
if pc = 46908 then
	inst <= x"C43C0010";
end if;
if pc = 46912 then
	inst <= x"C45C0014";
end if;
if pc = 46916 then
	inst <= x"C17DFFFC";
end if;
if pc = 46920 then
	inst <= x"00260000";
end if;
if pc = 46924 then
	inst <= x"03DC0020";
end if;
if pc = 46928 then
	inst <= x"037E000C";
end if;
if pc = 46932 then
	inst <= x"C57DFFFC";
end if;
if pc = 46936 then
	inst <= x"8200081C";
end if;
if pc = 46940 then
	inst <= x"07DC0020";
end if;
if pc = 46944 then
	inst <= x"005A0000";
end if;
if pc = 46948 then
	inst <= x"03BA0008";
end if;
if pc = 46952 then
	inst <= x"C4240004";
end if;
if pc = 46956 then
	inst <= x"C03C0014";
end if;
if pc = 46960 then
	inst <= x"C4240000";
end if;
if pc = 46964 then
	inst <= x"00240000";
end if;
if pc = 46968 then
	inst <= x"C05C000C";
end if;
if pc = 46972 then
	inst <= x"22640220";
end if;
if pc = 46976 then
	inst <= x"C09C0008";
end if;
if pc = 46980 then
	inst <= x"D4286000";
end if;
if pc = 46984 then
	inst <= x"06240001";
end if;
if pc = 46988 then
	inst <= x"8620B924";
end if;
if pc = 46992 then
	inst <= x"02400003";
end if;
if pc = 46996 then
	inst <= x"C83C0000";
end if;
if pc = 47000 then
	inst <= x"C43C0018";
end if;
if pc = 47004 then
	inst <= x"C17DFFFC";
end if;
if pc = 47008 then
	inst <= x"00240000";
end if;
if pc = 47012 then
	inst <= x"03DC0024";
end if;
if pc = 47016 then
	inst <= x"037E000C";
end if;
if pc = 47020 then
	inst <= x"C57DFFFC";
end if;
if pc = 47024 then
	inst <= x"8200081C";
end if;
if pc = 47028 then
	inst <= x"07DC0024";
end if;
if pc = 47032 then
	inst <= x"00420000";
end if;
if pc = 47036 then
	inst <= x"C03C0010";
end if;
if pc = 47040 then
	inst <= x"C0620000";
end if;
if pc = 47044 then
	inst <= x"C45C001C";
end if;
if pc = 47048 then
	inst <= x"C17DFFFC";
end if;
if pc = 47052 then
	inst <= x"00260000";
end if;
if pc = 47056 then
	inst <= x"03DC0028";
end if;
if pc = 47060 then
	inst <= x"037E000C";
end if;
if pc = 47064 then
	inst <= x"C57DFFFC";
end if;
if pc = 47068 then
	inst <= x"8200081C";
end if;
if pc = 47072 then
	inst <= x"07DC0028";
end if;
if pc = 47076 then
	inst <= x"005A0000";
end if;
if pc = 47080 then
	inst <= x"03BA0008";
end if;
if pc = 47084 then
	inst <= x"C4240004";
end if;
if pc = 47088 then
	inst <= x"C03C001C";
end if;
if pc = 47092 then
	inst <= x"C4240000";
end if;
if pc = 47096 then
	inst <= x"00240000";
end if;
if pc = 47100 then
	inst <= x"C05C0018";
end if;
if pc = 47104 then
	inst <= x"22640220";
end if;
if pc = 47108 then
	inst <= x"C09C0008";
end if;
if pc = 47112 then
	inst <= x"D4286000";
end if;
if pc = 47116 then
	inst <= x"06240001";
end if;
if pc = 47120 then
	inst <= x"8620B920";
end if;
if pc = 47124 then
	inst <= x"02400003";
end if;
if pc = 47128 then
	inst <= x"C83C0000";
end if;
if pc = 47132 then
	inst <= x"C43C0020";
end if;
if pc = 47136 then
	inst <= x"C17DFFFC";
end if;
if pc = 47140 then
	inst <= x"00240000";
end if;
if pc = 47144 then
	inst <= x"03DC002C";
end if;
if pc = 47148 then
	inst <= x"037E000C";
end if;
if pc = 47152 then
	inst <= x"C57DFFFC";
end if;
if pc = 47156 then
	inst <= x"8200081C";
end if;
if pc = 47160 then
	inst <= x"07DC002C";
end if;
if pc = 47164 then
	inst <= x"00420000";
end if;
if pc = 47168 then
	inst <= x"C03C0010";
end if;
if pc = 47172 then
	inst <= x"C0620000";
end if;
if pc = 47176 then
	inst <= x"C45C0024";
end if;
if pc = 47180 then
	inst <= x"C17DFFFC";
end if;
if pc = 47184 then
	inst <= x"00260000";
end if;
if pc = 47188 then
	inst <= x"03DC0030";
end if;
if pc = 47192 then
	inst <= x"037E000C";
end if;
if pc = 47196 then
	inst <= x"C57DFFFC";
end if;
if pc = 47200 then
	inst <= x"8200081C";
end if;
if pc = 47204 then
	inst <= x"07DC0030";
end if;
if pc = 47208 then
	inst <= x"005A0000";
end if;
if pc = 47212 then
	inst <= x"03BA0008";
end if;
if pc = 47216 then
	inst <= x"C4240004";
end if;
if pc = 47220 then
	inst <= x"C03C0024";
end if;
if pc = 47224 then
	inst <= x"C4240000";
end if;
if pc = 47228 then
	inst <= x"00240000";
end if;
if pc = 47232 then
	inst <= x"C05C0020";
end if;
if pc = 47236 then
	inst <= x"22640220";
end if;
if pc = 47240 then
	inst <= x"C09C0008";
end if;
if pc = 47244 then
	inst <= x"D4286000";
end if;
if pc = 47248 then
	inst <= x"06240001";
end if;
if pc = 47252 then
	inst <= x"8620B91C";
end if;
if pc = 47256 then
	inst <= x"02400003";
end if;
if pc = 47260 then
	inst <= x"C83C0000";
end if;
if pc = 47264 then
	inst <= x"C43C0028";
end if;
if pc = 47268 then
	inst <= x"C17DFFFC";
end if;
if pc = 47272 then
	inst <= x"00240000";
end if;
if pc = 47276 then
	inst <= x"03DC0034";
end if;
if pc = 47280 then
	inst <= x"037E000C";
end if;
if pc = 47284 then
	inst <= x"C57DFFFC";
end if;
if pc = 47288 then
	inst <= x"8200081C";
end if;
if pc = 47292 then
	inst <= x"07DC0034";
end if;
if pc = 47296 then
	inst <= x"00420000";
end if;
if pc = 47300 then
	inst <= x"C03C0010";
end if;
if pc = 47304 then
	inst <= x"C0220000";
end if;
if pc = 47308 then
	inst <= x"C45C002C";
end if;
if pc = 47312 then
	inst <= x"C17DFFFC";
end if;
if pc = 47316 then
	inst <= x"03DC0038";
end if;
if pc = 47320 then
	inst <= x"037E000C";
end if;
if pc = 47324 then
	inst <= x"C57DFFFC";
end if;
if pc = 47328 then
	inst <= x"8200081C";
end if;
if pc = 47332 then
	inst <= x"07DC0038";
end if;
if pc = 47336 then
	inst <= x"005A0000";
end if;
if pc = 47340 then
	inst <= x"03BA0008";
end if;
if pc = 47344 then
	inst <= x"C4240004";
end if;
if pc = 47348 then
	inst <= x"C03C002C";
end if;
if pc = 47352 then
	inst <= x"C4240000";
end if;
if pc = 47356 then
	inst <= x"00240000";
end if;
if pc = 47360 then
	inst <= x"C05C0028";
end if;
if pc = 47364 then
	inst <= x"22640220";
end if;
if pc = 47368 then
	inst <= x"C09C0008";
end if;
if pc = 47372 then
	inst <= x"D4286000";
end if;
if pc = 47376 then
	inst <= x"06440001";
end if;
if pc = 47380 then
	inst <= x"00280000";
end if;
if pc = 47384 then
	inst <= x"8200B6FC";
end if;
if pc = 47388 then
	inst <= x"C1FDFFFC";
end if;
if pc = 47392 then
	inst <= x"C1FDFFFC";
end if;
if pc = 47396 then
	inst <= x"C1FDFFFC";
end if;
if pc = 47400 then
	inst <= x"C1FDFFFC";
end if;
if pc = 47404 then
	inst <= x"8620BD0C";
end if;
if pc = 47408 then
	inst <= x"02400354";
end if;
if pc = 47412 then
	inst <= x"02600078";
end if;
if pc = 47416 then
	inst <= x"02800003";
end if;
if pc = 47420 then
	inst <= x"40200000";
end if;
if pc = 47424 then
	inst <= x"CC3C0000";
end if;
if pc = 47428 then
	inst <= x"C45C0008";
end if;
if pc = 47432 then
	inst <= x"C43C000C";
end if;
if pc = 47436 then
	inst <= x"C47C0010";
end if;
if pc = 47440 then
	inst <= x"C17DFFFC";
end if;
if pc = 47444 then
	inst <= x"00280000";
end if;
if pc = 47448 then
	inst <= x"03DC001C";
end if;
if pc = 47452 then
	inst <= x"037E000C";
end if;
if pc = 47456 then
	inst <= x"C57DFFFC";
end if;
if pc = 47460 then
	inst <= x"8200081C";
end if;
if pc = 47464 then
	inst <= x"07DC001C";
end if;
if pc = 47468 then
	inst <= x"00420000";
end if;
if pc = 47472 then
	inst <= x"022000C4";
end if;
if pc = 47476 then
	inst <= x"C0620000";
end if;
if pc = 47480 then
	inst <= x"C43C0014";
end if;
if pc = 47484 then
	inst <= x"C45C0018";
end if;
if pc = 47488 then
	inst <= x"C17DFFFC";
end if;
if pc = 47492 then
	inst <= x"00260000";
end if;
if pc = 47496 then
	inst <= x"03DC0024";
end if;
if pc = 47500 then
	inst <= x"037E000C";
end if;
if pc = 47504 then
	inst <= x"C57DFFFC";
end if;
if pc = 47508 then
	inst <= x"8200081C";
end if;
if pc = 47512 then
	inst <= x"07DC0024";
end if;
if pc = 47516 then
	inst <= x"005A0000";
end if;
if pc = 47520 then
	inst <= x"03BA0008";
end if;
if pc = 47524 then
	inst <= x"C4240004";
end if;
if pc = 47528 then
	inst <= x"C03C0018";
end if;
if pc = 47532 then
	inst <= x"C4240000";
end if;
if pc = 47536 then
	inst <= x"C03C0010";
end if;
if pc = 47540 then
	inst <= x"C17DFFFC";
end if;
if pc = 47544 then
	inst <= x"03DC0024";
end if;
if pc = 47548 then
	inst <= x"037E000C";
end if;
if pc = 47552 then
	inst <= x"C57DFFFC";
end if;
if pc = 47556 then
	inst <= x"8200081C";
end if;
if pc = 47560 then
	inst <= x"07DC0024";
end if;
if pc = 47564 then
	inst <= x"C05C000C";
end if;
if pc = 47568 then
	inst <= x"22640220";
end if;
if pc = 47572 then
	inst <= x"C09C0008";
end if;
if pc = 47576 then
	inst <= x"D4286000";
end if;
if pc = 47580 then
	inst <= x"02600003";
end if;
if pc = 47584 then
	inst <= x"C83C0000";
end if;
if pc = 47588 then
	inst <= x"C43C001C";
end if;
if pc = 47592 then
	inst <= x"C17DFFFC";
end if;
if pc = 47596 then
	inst <= x"00260000";
end if;
if pc = 47600 then
	inst <= x"03DC0028";
end if;
if pc = 47604 then
	inst <= x"037E000C";
end if;
if pc = 47608 then
	inst <= x"C57DFFFC";
end if;
if pc = 47612 then
	inst <= x"8200081C";
end if;
if pc = 47616 then
	inst <= x"07DC0028";
end if;
if pc = 47620 then
	inst <= x"00420000";
end if;
if pc = 47624 then
	inst <= x"C03C0014";
end if;
if pc = 47628 then
	inst <= x"C0620000";
end if;
if pc = 47632 then
	inst <= x"C45C0020";
end if;
if pc = 47636 then
	inst <= x"C17DFFFC";
end if;
if pc = 47640 then
	inst <= x"00260000";
end if;
if pc = 47644 then
	inst <= x"03DC002C";
end if;
if pc = 47648 then
	inst <= x"037E000C";
end if;
if pc = 47652 then
	inst <= x"C57DFFFC";
end if;
if pc = 47656 then
	inst <= x"8200081C";
end if;
if pc = 47660 then
	inst <= x"07DC002C";
end if;
if pc = 47664 then
	inst <= x"005A0000";
end if;
if pc = 47668 then
	inst <= x"03BA0008";
end if;
if pc = 47672 then
	inst <= x"C4240004";
end if;
if pc = 47676 then
	inst <= x"C03C0020";
end if;
if pc = 47680 then
	inst <= x"C4240000";
end if;
if pc = 47684 then
	inst <= x"00240000";
end if;
if pc = 47688 then
	inst <= x"C05C001C";
end if;
if pc = 47692 then
	inst <= x"C42401D8";
end if;
if pc = 47696 then
	inst <= x"02200003";
end if;
if pc = 47700 then
	inst <= x"C83C0000";
end if;
if pc = 47704 then
	inst <= x"C17DFFFC";
end if;
if pc = 47708 then
	inst <= x"03DC002C";
end if;
if pc = 47712 then
	inst <= x"037E000C";
end if;
if pc = 47716 then
	inst <= x"C57DFFFC";
end if;
if pc = 47720 then
	inst <= x"8200081C";
end if;
if pc = 47724 then
	inst <= x"07DC002C";
end if;
if pc = 47728 then
	inst <= x"00420000";
end if;
if pc = 47732 then
	inst <= x"C03C0014";
end if;
if pc = 47736 then
	inst <= x"C0620000";
end if;
if pc = 47740 then
	inst <= x"C45C0024";
end if;
if pc = 47744 then
	inst <= x"C17DFFFC";
end if;
if pc = 47748 then
	inst <= x"00260000";
end if;
if pc = 47752 then
	inst <= x"03DC0030";
end if;
if pc = 47756 then
	inst <= x"037E000C";
end if;
if pc = 47760 then
	inst <= x"C57DFFFC";
end if;
if pc = 47764 then
	inst <= x"8200081C";
end if;
if pc = 47768 then
	inst <= x"07DC0030";
end if;
if pc = 47772 then
	inst <= x"005A0000";
end if;
if pc = 47776 then
	inst <= x"03BA0008";
end if;
if pc = 47780 then
	inst <= x"C4240004";
end if;
if pc = 47784 then
	inst <= x"C03C0024";
end if;
if pc = 47788 then
	inst <= x"C4240000";
end if;
if pc = 47792 then
	inst <= x"00240000";
end if;
if pc = 47796 then
	inst <= x"C05C001C";
end if;
if pc = 47800 then
	inst <= x"C42401D4";
end if;
if pc = 47804 then
	inst <= x"02200003";
end if;
if pc = 47808 then
	inst <= x"C83C0000";
end if;
if pc = 47812 then
	inst <= x"C17DFFFC";
end if;
if pc = 47816 then
	inst <= x"03DC0030";
end if;
if pc = 47820 then
	inst <= x"037E000C";
end if;
if pc = 47824 then
	inst <= x"C57DFFFC";
end if;
if pc = 47828 then
	inst <= x"8200081C";
end if;
if pc = 47832 then
	inst <= x"07DC0030";
end if;
if pc = 47836 then
	inst <= x"00420000";
end if;
if pc = 47840 then
	inst <= x"C03C0014";
end if;
if pc = 47844 then
	inst <= x"C0620000";
end if;
if pc = 47848 then
	inst <= x"C45C0028";
end if;
if pc = 47852 then
	inst <= x"C17DFFFC";
end if;
if pc = 47856 then
	inst <= x"00260000";
end if;
if pc = 47860 then
	inst <= x"03DC0034";
end if;
if pc = 47864 then
	inst <= x"037E000C";
end if;
if pc = 47868 then
	inst <= x"C57DFFFC";
end if;
if pc = 47872 then
	inst <= x"8200081C";
end if;
if pc = 47876 then
	inst <= x"07DC0034";
end if;
if pc = 47880 then
	inst <= x"005A0000";
end if;
if pc = 47884 then
	inst <= x"03BA0008";
end if;
if pc = 47888 then
	inst <= x"C4240004";
end if;
if pc = 47892 then
	inst <= x"C03C0028";
end if;
if pc = 47896 then
	inst <= x"C4240000";
end if;
if pc = 47900 then
	inst <= x"00240000";
end if;
if pc = 47904 then
	inst <= x"C05C001C";
end if;
if pc = 47908 then
	inst <= x"C42401D0";
end if;
if pc = 47912 then
	inst <= x"02200073";
end if;
if pc = 47916 then
	inst <= x"C17DFFFC";
end if;
if pc = 47920 then
	inst <= x"01240000";
end if;
if pc = 47924 then
	inst <= x"00420000";
end if;
if pc = 47928 then
	inst <= x"00320000";
end if;
if pc = 47932 then
	inst <= x"03DC0034";
end if;
if pc = 47936 then
	inst <= x"037E000C";
end if;
if pc = 47940 then
	inst <= x"C57DFFFC";
end if;
if pc = 47944 then
	inst <= x"8200B6FC";
end if;
if pc = 47948 then
	inst <= x"07DC0034";
end if;
if pc = 47952 then
	inst <= x"C03C000C";
end if;
if pc = 47956 then
	inst <= x"06220001";
end if;
if pc = 47960 then
	inst <= x"8620BD08";
end if;
if pc = 47964 then
	inst <= x"02400078";
end if;
if pc = 47968 then
	inst <= x"02600003";
end if;
if pc = 47972 then
	inst <= x"C83C0000";
end if;
if pc = 47976 then
	inst <= x"C43C002C";
end if;
if pc = 47980 then
	inst <= x"C45C0030";
end if;
if pc = 47984 then
	inst <= x"C17DFFFC";
end if;
if pc = 47988 then
	inst <= x"00260000";
end if;
if pc = 47992 then
	inst <= x"03DC003C";
end if;
if pc = 47996 then
	inst <= x"037E000C";
end if;
if pc = 48000 then
	inst <= x"C57DFFFC";
end if;
if pc = 48004 then
	inst <= x"8200081C";
end if;
if pc = 48008 then
	inst <= x"07DC003C";
end if;
if pc = 48012 then
	inst <= x"00420000";
end if;
if pc = 48016 then
	inst <= x"C03C0014";
end if;
if pc = 48020 then
	inst <= x"C0620000";
end if;
if pc = 48024 then
	inst <= x"C45C0034";
end if;
if pc = 48028 then
	inst <= x"C17DFFFC";
end if;
if pc = 48032 then
	inst <= x"00260000";
end if;
if pc = 48036 then
	inst <= x"03DC0040";
end if;
if pc = 48040 then
	inst <= x"037E000C";
end if;
if pc = 48044 then
	inst <= x"C57DFFFC";
end if;
if pc = 48048 then
	inst <= x"8200081C";
end if;
if pc = 48052 then
	inst <= x"07DC0040";
end if;
if pc = 48056 then
	inst <= x"005A0000";
end if;
if pc = 48060 then
	inst <= x"03BA0008";
end if;
if pc = 48064 then
	inst <= x"C4240004";
end if;
if pc = 48068 then
	inst <= x"C03C0034";
end if;
if pc = 48072 then
	inst <= x"C4240000";
end if;
if pc = 48076 then
	inst <= x"C03C0030";
end if;
if pc = 48080 then
	inst <= x"C17DFFFC";
end if;
if pc = 48084 then
	inst <= x"03DC0040";
end if;
if pc = 48088 then
	inst <= x"037E000C";
end if;
if pc = 48092 then
	inst <= x"C57DFFFC";
end if;
if pc = 48096 then
	inst <= x"8200081C";
end if;
if pc = 48100 then
	inst <= x"07DC0040";
end if;
if pc = 48104 then
	inst <= x"C05C002C";
end if;
if pc = 48108 then
	inst <= x"22640220";
end if;
if pc = 48112 then
	inst <= x"C09C0008";
end if;
if pc = 48116 then
	inst <= x"D4286000";
end if;
if pc = 48120 then
	inst <= x"02600003";
end if;
if pc = 48124 then
	inst <= x"C83C0000";
end if;
if pc = 48128 then
	inst <= x"C43C0038";
end if;
if pc = 48132 then
	inst <= x"C17DFFFC";
end if;
if pc = 48136 then
	inst <= x"00260000";
end if;
if pc = 48140 then
	inst <= x"03DC0044";
end if;
if pc = 48144 then
	inst <= x"037E000C";
end if;
if pc = 48148 then
	inst <= x"C57DFFFC";
end if;
if pc = 48152 then
	inst <= x"8200081C";
end if;
if pc = 48156 then
	inst <= x"07DC0044";
end if;
if pc = 48160 then
	inst <= x"00420000";
end if;
if pc = 48164 then
	inst <= x"C03C0014";
end if;
if pc = 48168 then
	inst <= x"C0620000";
end if;
if pc = 48172 then
	inst <= x"C45C003C";
end if;
if pc = 48176 then
	inst <= x"C17DFFFC";
end if;
if pc = 48180 then
	inst <= x"00260000";
end if;
if pc = 48184 then
	inst <= x"03DC0048";
end if;
if pc = 48188 then
	inst <= x"037E000C";
end if;
if pc = 48192 then
	inst <= x"C57DFFFC";
end if;
if pc = 48196 then
	inst <= x"8200081C";
end if;
if pc = 48200 then
	inst <= x"07DC0048";
end if;
if pc = 48204 then
	inst <= x"005A0000";
end if;
if pc = 48208 then
	inst <= x"03BA0008";
end if;
if pc = 48212 then
	inst <= x"C4240004";
end if;
if pc = 48216 then
	inst <= x"C03C003C";
end if;
if pc = 48220 then
	inst <= x"C4240000";
end if;
if pc = 48224 then
	inst <= x"00240000";
end if;
if pc = 48228 then
	inst <= x"C05C0038";
end if;
if pc = 48232 then
	inst <= x"C42401D8";
end if;
if pc = 48236 then
	inst <= x"02200003";
end if;
if pc = 48240 then
	inst <= x"C83C0000";
end if;
if pc = 48244 then
	inst <= x"C17DFFFC";
end if;
if pc = 48248 then
	inst <= x"03DC0048";
end if;
if pc = 48252 then
	inst <= x"037E000C";
end if;
if pc = 48256 then
	inst <= x"C57DFFFC";
end if;
if pc = 48260 then
	inst <= x"8200081C";
end if;
if pc = 48264 then
	inst <= x"07DC0048";
end if;
if pc = 48268 then
	inst <= x"00420000";
end if;
if pc = 48272 then
	inst <= x"C03C0014";
end if;
if pc = 48276 then
	inst <= x"C0220000";
end if;
if pc = 48280 then
	inst <= x"C45C0040";
end if;
if pc = 48284 then
	inst <= x"C17DFFFC";
end if;
if pc = 48288 then
	inst <= x"03DC004C";
end if;
if pc = 48292 then
	inst <= x"037E000C";
end if;
if pc = 48296 then
	inst <= x"C57DFFFC";
end if;
if pc = 48300 then
	inst <= x"8200081C";
end if;
if pc = 48304 then
	inst <= x"07DC004C";
end if;
if pc = 48308 then
	inst <= x"005A0000";
end if;
if pc = 48312 then
	inst <= x"03BA0008";
end if;
if pc = 48316 then
	inst <= x"C4240004";
end if;
if pc = 48320 then
	inst <= x"C03C0040";
end if;
if pc = 48324 then
	inst <= x"C4240000";
end if;
if pc = 48328 then
	inst <= x"00240000";
end if;
if pc = 48332 then
	inst <= x"C05C0038";
end if;
if pc = 48336 then
	inst <= x"C42401D4";
end if;
if pc = 48340 then
	inst <= x"02200074";
end if;
if pc = 48344 then
	inst <= x"C17DFFFC";
end if;
if pc = 48348 then
	inst <= x"01240000";
end if;
if pc = 48352 then
	inst <= x"00420000";
end if;
if pc = 48356 then
	inst <= x"00320000";
end if;
if pc = 48360 then
	inst <= x"03DC004C";
end if;
if pc = 48364 then
	inst <= x"037E000C";
end if;
if pc = 48368 then
	inst <= x"C57DFFFC";
end if;
if pc = 48372 then
	inst <= x"8200B6FC";
end if;
if pc = 48376 then
	inst <= x"07DC004C";
end if;
if pc = 48380 then
	inst <= x"C03C002C";
end if;
if pc = 48384 then
	inst <= x"06220001";
end if;
if pc = 48388 then
	inst <= x"8200B92C";
end if;
if pc = 48392 then
	inst <= x"C1FDFFFC";
end if;
if pc = 48396 then
	inst <= x"C1FDFFFC";
end if;
if pc = 48400 then
	inst <= x"8640C710";
end if;
if pc = 48404 then
	inst <= x"22640220";
end if;
if pc = 48408 then
	inst <= x"D0626000";
end if;
if pc = 48412 then
	inst <= x"028000C4";
end if;
if pc = 48416 then
	inst <= x"C0A80000";
end if;
if pc = 48420 then
	inst <= x"06AA0001";
end if;
if pc = 48424 then
	inst <= x"C49C0000";
end if;
if pc = 48428 then
	inst <= x"C43C0004";
end if;
if pc = 48432 then
	inst <= x"C45C0008";
end if;
if pc = 48436 then
	inst <= x"86A0BF18";
end if;
if pc = 48440 then
	inst <= x"02C000C8";
end if;
if pc = 48444 then
	inst <= x"22EA0220";
end if;
if pc = 48448 then
	inst <= x"D0ECE000";
end if;
if pc = 48452 then
	inst <= x"C1060004";
end if;
if pc = 48456 then
	inst <= x"C1260000";
end if;
if pc = 48460 then
	inst <= x"C14E0004";
end if;
if pc = 48464 then
	inst <= x"02800001";
end if;
if pc = 48468 then
	inst <= x"C47C000C";
end if;
if pc = 48472 then
	inst <= x"C4DC0010";
end if;
if pc = 48476 then
	inst <= x"8348BDE0";
end if;
if pc = 48480 then
	inst <= x"02800002";
end if;
if pc = 48484 then
	inst <= x"8348BDA4";
end if;
if pc = 48488 then
	inst <= x"C51C0014";
end if;
if pc = 48492 then
	inst <= x"C4BC0018";
end if;
if pc = 48496 then
	inst <= x"C17DFFFC";
end if;
if pc = 48500 then
	inst <= x"004E0000";
end if;
if pc = 48504 then
	inst <= x"00320000";
end if;
if pc = 48508 then
	inst <= x"03DC0024";
end if;
if pc = 48512 then
	inst <= x"037E000C";
end if;
if pc = 48516 then
	inst <= x"C57DFFFC";
end if;
if pc = 48520 then
	inst <= x"8200400C";
end if;
if pc = 48524 then
	inst <= x"07DC0024";
end if;
if pc = 48528 then
	inst <= x"C05C0018";
end if;
if pc = 48532 then
	inst <= x"22640220";
end if;
if pc = 48536 then
	inst <= x"C09C0014";
end if;
if pc = 48540 then
	inst <= x"D4286000";
end if;
if pc = 48544 then
	inst <= x"8200BDDC";
end if;
if pc = 48548 then
	inst <= x"C51C0014";
end if;
if pc = 48552 then
	inst <= x"C4BC0018";
end if;
if pc = 48556 then
	inst <= x"C17DFFFC";
end if;
if pc = 48560 then
	inst <= x"004E0000";
end if;
if pc = 48564 then
	inst <= x"00320000";
end if;
if pc = 48568 then
	inst <= x"03DC0024";
end if;
if pc = 48572 then
	inst <= x"037E000C";
end if;
if pc = 48576 then
	inst <= x"C57DFFFC";
end if;
if pc = 48580 then
	inst <= x"82003E98";
end if;
if pc = 48584 then
	inst <= x"07DC0024";
end if;
if pc = 48588 then
	inst <= x"C05C0018";
end if;
if pc = 48592 then
	inst <= x"22640220";
end if;
if pc = 48596 then
	inst <= x"C09C0014";
end if;
if pc = 48600 then
	inst <= x"D4286000";
end if;
if pc = 48604 then
	inst <= x"8200BE18";
end if;
if pc = 48608 then
	inst <= x"C51C0014";
end if;
if pc = 48612 then
	inst <= x"C4BC0018";
end if;
if pc = 48616 then
	inst <= x"C17DFFFC";
end if;
if pc = 48620 then
	inst <= x"004E0000";
end if;
if pc = 48624 then
	inst <= x"00320000";
end if;
if pc = 48628 then
	inst <= x"03DC0024";
end if;
if pc = 48632 then
	inst <= x"037E000C";
end if;
if pc = 48636 then
	inst <= x"C57DFFFC";
end if;
if pc = 48640 then
	inst <= x"82003CC4";
end if;
if pc = 48644 then
	inst <= x"07DC0024";
end if;
if pc = 48648 then
	inst <= x"C05C0018";
end if;
if pc = 48652 then
	inst <= x"22640220";
end if;
if pc = 48656 then
	inst <= x"C09C0014";
end if;
if pc = 48660 then
	inst <= x"D4286000";
end if;
if pc = 48664 then
	inst <= x"06240001";
end if;
if pc = 48668 then
	inst <= x"8620BF14";
end if;
if pc = 48672 then
	inst <= x"22420220";
end if;
if pc = 48676 then
	inst <= x"C07C0010";
end if;
if pc = 48680 then
	inst <= x"D0464000";
end if;
if pc = 48684 then
	inst <= x"C07C000C";
end if;
if pc = 48688 then
	inst <= x"C0860004";
end if;
if pc = 48692 then
	inst <= x"C0A60000";
end if;
if pc = 48696 then
	inst <= x"C0C40004";
end if;
if pc = 48700 then
	inst <= x"02E00001";
end if;
if pc = 48704 then
	inst <= x"82CEBEBC";
end if;
if pc = 48708 then
	inst <= x"02E00002";
end if;
if pc = 48712 then
	inst <= x"82CEBE84";
end if;
if pc = 48716 then
	inst <= x"C49C001C";
end if;
if pc = 48720 then
	inst <= x"C43C0020";
end if;
if pc = 48724 then
	inst <= x"C17DFFFC";
end if;
if pc = 48728 then
	inst <= x"002A0000";
end if;
if pc = 48732 then
	inst <= x"03DC002C";
end if;
if pc = 48736 then
	inst <= x"037E000C";
end if;
if pc = 48740 then
	inst <= x"C57DFFFC";
end if;
if pc = 48744 then
	inst <= x"8200400C";
end if;
if pc = 48748 then
	inst <= x"07DC002C";
end if;
if pc = 48752 then
	inst <= x"C05C0020";
end if;
if pc = 48756 then
	inst <= x"22640220";
end if;
if pc = 48760 then
	inst <= x"C09C001C";
end if;
if pc = 48764 then
	inst <= x"D4286000";
end if;
if pc = 48768 then
	inst <= x"8200BEB8";
end if;
if pc = 48772 then
	inst <= x"C49C001C";
end if;
if pc = 48776 then
	inst <= x"C43C0020";
end if;
if pc = 48780 then
	inst <= x"C17DFFFC";
end if;
if pc = 48784 then
	inst <= x"002A0000";
end if;
if pc = 48788 then
	inst <= x"03DC002C";
end if;
if pc = 48792 then
	inst <= x"037E000C";
end if;
if pc = 48796 then
	inst <= x"C57DFFFC";
end if;
if pc = 48800 then
	inst <= x"82003E98";
end if;
if pc = 48804 then
	inst <= x"07DC002C";
end if;
if pc = 48808 then
	inst <= x"C05C0020";
end if;
if pc = 48812 then
	inst <= x"22640220";
end if;
if pc = 48816 then
	inst <= x"C09C001C";
end if;
if pc = 48820 then
	inst <= x"D4286000";
end if;
if pc = 48824 then
	inst <= x"8200BEF0";
end if;
if pc = 48828 then
	inst <= x"C49C001C";
end if;
if pc = 48832 then
	inst <= x"C43C0020";
end if;
if pc = 48836 then
	inst <= x"C17DFFFC";
end if;
if pc = 48840 then
	inst <= x"002A0000";
end if;
if pc = 48844 then
	inst <= x"03DC002C";
end if;
if pc = 48848 then
	inst <= x"037E000C";
end if;
if pc = 48852 then
	inst <= x"C57DFFFC";
end if;
if pc = 48856 then
	inst <= x"82003CC4";
end if;
if pc = 48860 then
	inst <= x"07DC002C";
end if;
if pc = 48864 then
	inst <= x"C05C0020";
end if;
if pc = 48868 then
	inst <= x"22640220";
end if;
if pc = 48872 then
	inst <= x"C09C001C";
end if;
if pc = 48876 then
	inst <= x"D4286000";
end if;
if pc = 48880 then
	inst <= x"06440001";
end if;
if pc = 48884 then
	inst <= x"C03C000C";
end if;
if pc = 48888 then
	inst <= x"C17DFFFC";
end if;
if pc = 48892 then
	inst <= x"03DC002C";
end if;
if pc = 48896 then
	inst <= x"037E000C";
end if;
if pc = 48900 then
	inst <= x"C57DFFFC";
end if;
if pc = 48904 then
	inst <= x"820042A4";
end if;
if pc = 48908 then
	inst <= x"07DC002C";
end if;
if pc = 48912 then
	inst <= x"8200BF14";
end if;
if pc = 48916 then
	inst <= x"8200BF18";
end if;
if pc = 48920 then
	inst <= x"C03C0008";
end if;
if pc = 48924 then
	inst <= x"06220001";
end if;
if pc = 48928 then
	inst <= x"8620C70C";
end if;
if pc = 48932 then
	inst <= x"22420220";
end if;
if pc = 48936 then
	inst <= x"C07C0004";
end if;
if pc = 48940 then
	inst <= x"D0464000";
end if;
if pc = 48944 then
	inst <= x"C09C0000";
end if;
if pc = 48948 then
	inst <= x"C0A80000";
end if;
if pc = 48952 then
	inst <= x"06AA0001";
end if;
if pc = 48956 then
	inst <= x"C43C0024";
end if;
if pc = 48960 then
	inst <= x"86A0C200";
end if;
if pc = 48964 then
	inst <= x"02C000C8";
end if;
if pc = 48968 then
	inst <= x"22EA0220";
end if;
if pc = 48972 then
	inst <= x"D0ECE000";
end if;
if pc = 48976 then
	inst <= x"C1040004";
end if;
if pc = 48980 then
	inst <= x"C1240000";
end if;
if pc = 48984 then
	inst <= x"C14E0004";
end if;
if pc = 48988 then
	inst <= x"02800001";
end if;
if pc = 48992 then
	inst <= x"C45C0028";
end if;
if pc = 48996 then
	inst <= x"C4DC002C";
end if;
if pc = 49000 then
	inst <= x"8348BFEC";
end if;
if pc = 49004 then
	inst <= x"02800002";
end if;
if pc = 49008 then
	inst <= x"8348BFB0";
end if;
if pc = 49012 then
	inst <= x"C51C0030";
end if;
if pc = 49016 then
	inst <= x"C4BC0034";
end if;
if pc = 49020 then
	inst <= x"C17DFFFC";
end if;
if pc = 49024 then
	inst <= x"004E0000";
end if;
if pc = 49028 then
	inst <= x"00320000";
end if;
if pc = 49032 then
	inst <= x"03DC0040";
end if;
if pc = 49036 then
	inst <= x"037E000C";
end if;
if pc = 49040 then
	inst <= x"C57DFFFC";
end if;
if pc = 49044 then
	inst <= x"8200400C";
end if;
if pc = 49048 then
	inst <= x"07DC0040";
end if;
if pc = 49052 then
	inst <= x"C05C0034";
end if;
if pc = 49056 then
	inst <= x"22640220";
end if;
if pc = 49060 then
	inst <= x"C09C0030";
end if;
if pc = 49064 then
	inst <= x"D4286000";
end if;
if pc = 49068 then
	inst <= x"8200BFE8";
end if;
if pc = 49072 then
	inst <= x"C51C0030";
end if;
if pc = 49076 then
	inst <= x"C4BC0034";
end if;
if pc = 49080 then
	inst <= x"C17DFFFC";
end if;
if pc = 49084 then
	inst <= x"004E0000";
end if;
if pc = 49088 then
	inst <= x"00320000";
end if;
if pc = 49092 then
	inst <= x"03DC0040";
end if;
if pc = 49096 then
	inst <= x"037E000C";
end if;
if pc = 49100 then
	inst <= x"C57DFFFC";
end if;
if pc = 49104 then
	inst <= x"82003E98";
end if;
if pc = 49108 then
	inst <= x"07DC0040";
end if;
if pc = 49112 then
	inst <= x"C05C0034";
end if;
if pc = 49116 then
	inst <= x"22640220";
end if;
if pc = 49120 then
	inst <= x"C09C0030";
end if;
if pc = 49124 then
	inst <= x"D4286000";
end if;
if pc = 49128 then
	inst <= x"8200C024";
end if;
if pc = 49132 then
	inst <= x"C51C0030";
end if;
if pc = 49136 then
	inst <= x"C4BC0034";
end if;
if pc = 49140 then
	inst <= x"C17DFFFC";
end if;
if pc = 49144 then
	inst <= x"004E0000";
end if;
if pc = 49148 then
	inst <= x"00320000";
end if;
if pc = 49152 then
	inst <= x"03DC0040";
end if;
if pc = 49156 then
	inst <= x"037E000C";
end if;
if pc = 49160 then
	inst <= x"C57DFFFC";
end if;
if pc = 49164 then
	inst <= x"82003CC4";
end if;
if pc = 49168 then
	inst <= x"07DC0040";
end if;
if pc = 49172 then
	inst <= x"C05C0034";
end if;
if pc = 49176 then
	inst <= x"22640220";
end if;
if pc = 49180 then
	inst <= x"C09C0030";
end if;
if pc = 49184 then
	inst <= x"D4286000";
end if;
if pc = 49188 then
	inst <= x"06240001";
end if;
if pc = 49192 then
	inst <= x"8620C1FC";
end if;
if pc = 49196 then
	inst <= x"22420220";
end if;
if pc = 49200 then
	inst <= x"C07C002C";
end if;
if pc = 49204 then
	inst <= x"D0464000";
end if;
if pc = 49208 then
	inst <= x"C09C0028";
end if;
if pc = 49212 then
	inst <= x"C0A80004";
end if;
if pc = 49216 then
	inst <= x"C0C80000";
end if;
if pc = 49220 then
	inst <= x"C0E40004";
end if;
if pc = 49224 then
	inst <= x"03000001";
end if;
if pc = 49228 then
	inst <= x"82F0C0C8";
end if;
if pc = 49232 then
	inst <= x"03000002";
end if;
if pc = 49236 then
	inst <= x"82F0C090";
end if;
if pc = 49240 then
	inst <= x"C4BC0038";
end if;
if pc = 49244 then
	inst <= x"C43C003C";
end if;
if pc = 49248 then
	inst <= x"C17DFFFC";
end if;
if pc = 49252 then
	inst <= x"002C0000";
end if;
if pc = 49256 then
	inst <= x"03DC0048";
end if;
if pc = 49260 then
	inst <= x"037E000C";
end if;
if pc = 49264 then
	inst <= x"C57DFFFC";
end if;
if pc = 49268 then
	inst <= x"8200400C";
end if;
if pc = 49272 then
	inst <= x"07DC0048";
end if;
if pc = 49276 then
	inst <= x"C05C003C";
end if;
if pc = 49280 then
	inst <= x"22640220";
end if;
if pc = 49284 then
	inst <= x"C09C0038";
end if;
if pc = 49288 then
	inst <= x"D4286000";
end if;
if pc = 49292 then
	inst <= x"8200C0C4";
end if;
if pc = 49296 then
	inst <= x"C4BC0038";
end if;
if pc = 49300 then
	inst <= x"C43C003C";
end if;
if pc = 49304 then
	inst <= x"C17DFFFC";
end if;
if pc = 49308 then
	inst <= x"002C0000";
end if;
if pc = 49312 then
	inst <= x"03DC0048";
end if;
if pc = 49316 then
	inst <= x"037E000C";
end if;
if pc = 49320 then
	inst <= x"C57DFFFC";
end if;
if pc = 49324 then
	inst <= x"82003E98";
end if;
if pc = 49328 then
	inst <= x"07DC0048";
end if;
if pc = 49332 then
	inst <= x"C05C003C";
end if;
if pc = 49336 then
	inst <= x"22640220";
end if;
if pc = 49340 then
	inst <= x"C09C0038";
end if;
if pc = 49344 then
	inst <= x"D4286000";
end if;
if pc = 49348 then
	inst <= x"8200C0FC";
end if;
if pc = 49352 then
	inst <= x"C4BC0038";
end if;
if pc = 49356 then
	inst <= x"C43C003C";
end if;
if pc = 49360 then
	inst <= x"C17DFFFC";
end if;
if pc = 49364 then
	inst <= x"002C0000";
end if;
if pc = 49368 then
	inst <= x"03DC0048";
end if;
if pc = 49372 then
	inst <= x"037E000C";
end if;
if pc = 49376 then
	inst <= x"C57DFFFC";
end if;
if pc = 49380 then
	inst <= x"82003CC4";
end if;
if pc = 49384 then
	inst <= x"07DC0048";
end if;
if pc = 49388 then
	inst <= x"C05C003C";
end if;
if pc = 49392 then
	inst <= x"22640220";
end if;
if pc = 49396 then
	inst <= x"C09C0038";
end if;
if pc = 49400 then
	inst <= x"D4286000";
end if;
if pc = 49404 then
	inst <= x"06240001";
end if;
if pc = 49408 then
	inst <= x"8620C1F8";
end if;
if pc = 49412 then
	inst <= x"22420220";
end if;
if pc = 49416 then
	inst <= x"C07C002C";
end if;
if pc = 49420 then
	inst <= x"D0464000";
end if;
if pc = 49424 then
	inst <= x"C07C0028";
end if;
if pc = 49428 then
	inst <= x"C0860004";
end if;
if pc = 49432 then
	inst <= x"C0A60000";
end if;
if pc = 49436 then
	inst <= x"C0C40004";
end if;
if pc = 49440 then
	inst <= x"02E00001";
end if;
if pc = 49444 then
	inst <= x"82CEC1A0";
end if;
if pc = 49448 then
	inst <= x"02E00002";
end if;
if pc = 49452 then
	inst <= x"82CEC168";
end if;
if pc = 49456 then
	inst <= x"C49C0040";
end if;
if pc = 49460 then
	inst <= x"C43C0044";
end if;
if pc = 49464 then
	inst <= x"C17DFFFC";
end if;
if pc = 49468 then
	inst <= x"002A0000";
end if;
if pc = 49472 then
	inst <= x"03DC0050";
end if;
if pc = 49476 then
	inst <= x"037E000C";
end if;
if pc = 49480 then
	inst <= x"C57DFFFC";
end if;
if pc = 49484 then
	inst <= x"8200400C";
end if;
if pc = 49488 then
	inst <= x"07DC0050";
end if;
if pc = 49492 then
	inst <= x"C05C0044";
end if;
if pc = 49496 then
	inst <= x"22640220";
end if;
if pc = 49500 then
	inst <= x"C09C0040";
end if;
if pc = 49504 then
	inst <= x"D4286000";
end if;
if pc = 49508 then
	inst <= x"8200C19C";
end if;
if pc = 49512 then
	inst <= x"C49C0040";
end if;
if pc = 49516 then
	inst <= x"C43C0044";
end if;
if pc = 49520 then
	inst <= x"C17DFFFC";
end if;
if pc = 49524 then
	inst <= x"002A0000";
end if;
if pc = 49528 then
	inst <= x"03DC0050";
end if;
if pc = 49532 then
	inst <= x"037E000C";
end if;
if pc = 49536 then
	inst <= x"C57DFFFC";
end if;
if pc = 49540 then
	inst <= x"82003E98";
end if;
if pc = 49544 then
	inst <= x"07DC0050";
end if;
if pc = 49548 then
	inst <= x"C05C0044";
end if;
if pc = 49552 then
	inst <= x"22640220";
end if;
if pc = 49556 then
	inst <= x"C09C0040";
end if;
if pc = 49560 then
	inst <= x"D4286000";
end if;
if pc = 49564 then
	inst <= x"8200C1D4";
end if;
if pc = 49568 then
	inst <= x"C49C0040";
end if;
if pc = 49572 then
	inst <= x"C43C0044";
end if;
if pc = 49576 then
	inst <= x"C17DFFFC";
end if;
if pc = 49580 then
	inst <= x"002A0000";
end if;
if pc = 49584 then
	inst <= x"03DC0050";
end if;
if pc = 49588 then
	inst <= x"037E000C";
end if;
if pc = 49592 then
	inst <= x"C57DFFFC";
end if;
if pc = 49596 then
	inst <= x"82003CC4";
end if;
if pc = 49600 then
	inst <= x"07DC0050";
end if;
if pc = 49604 then
	inst <= x"C05C0044";
end if;
if pc = 49608 then
	inst <= x"22640220";
end if;
if pc = 49612 then
	inst <= x"C09C0040";
end if;
if pc = 49616 then
	inst <= x"D4286000";
end if;
if pc = 49620 then
	inst <= x"06440001";
end if;
if pc = 49624 then
	inst <= x"C03C0028";
end if;
if pc = 49628 then
	inst <= x"C17DFFFC";
end if;
if pc = 49632 then
	inst <= x"03DC0050";
end if;
if pc = 49636 then
	inst <= x"037E000C";
end if;
if pc = 49640 then
	inst <= x"C57DFFFC";
end if;
if pc = 49644 then
	inst <= x"820042A4";
end if;
if pc = 49648 then
	inst <= x"07DC0050";
end if;
if pc = 49652 then
	inst <= x"8200C1F8";
end if;
if pc = 49656 then
	inst <= x"8200C1FC";
end if;
if pc = 49660 then
	inst <= x"8200C200";
end if;
if pc = 49664 then
	inst <= x"C03C0024";
end if;
if pc = 49668 then
	inst <= x"06220001";
end if;
if pc = 49672 then
	inst <= x"8620C708";
end if;
if pc = 49676 then
	inst <= x"22420220";
end if;
if pc = 49680 then
	inst <= x"C07C0004";
end if;
if pc = 49684 then
	inst <= x"D0464000";
end if;
if pc = 49688 then
	inst <= x"C09C0000";
end if;
if pc = 49692 then
	inst <= x"C0A80000";
end if;
if pc = 49696 then
	inst <= x"06AA0001";
end if;
if pc = 49700 then
	inst <= x"C43C0048";
end if;
if pc = 49704 then
	inst <= x"86A0C40C";
end if;
if pc = 49708 then
	inst <= x"02C000C8";
end if;
if pc = 49712 then
	inst <= x"22EA0220";
end if;
if pc = 49716 then
	inst <= x"D0ECE000";
end if;
if pc = 49720 then
	inst <= x"C1040004";
end if;
if pc = 49724 then
	inst <= x"C1240000";
end if;
if pc = 49728 then
	inst <= x"C14E0004";
end if;
if pc = 49732 then
	inst <= x"02800001";
end if;
if pc = 49736 then
	inst <= x"C45C004C";
end if;
if pc = 49740 then
	inst <= x"C4DC0050";
end if;
if pc = 49744 then
	inst <= x"8348C2D4";
end if;
if pc = 49748 then
	inst <= x"02800002";
end if;
if pc = 49752 then
	inst <= x"8348C298";
end if;
if pc = 49756 then
	inst <= x"C51C0054";
end if;
if pc = 49760 then
	inst <= x"C4BC0058";
end if;
if pc = 49764 then
	inst <= x"C17DFFFC";
end if;
if pc = 49768 then
	inst <= x"004E0000";
end if;
if pc = 49772 then
	inst <= x"00320000";
end if;
if pc = 49776 then
	inst <= x"03DC0064";
end if;
if pc = 49780 then
	inst <= x"037E000C";
end if;
if pc = 49784 then
	inst <= x"C57DFFFC";
end if;
if pc = 49788 then
	inst <= x"8200400C";
end if;
if pc = 49792 then
	inst <= x"07DC0064";
end if;
if pc = 49796 then
	inst <= x"C05C0058";
end if;
if pc = 49800 then
	inst <= x"22640220";
end if;
if pc = 49804 then
	inst <= x"C09C0054";
end if;
if pc = 49808 then
	inst <= x"D4286000";
end if;
if pc = 49812 then
	inst <= x"8200C2D0";
end if;
if pc = 49816 then
	inst <= x"C51C0054";
end if;
if pc = 49820 then
	inst <= x"C4BC0058";
end if;
if pc = 49824 then
	inst <= x"C17DFFFC";
end if;
if pc = 49828 then
	inst <= x"004E0000";
end if;
if pc = 49832 then
	inst <= x"00320000";
end if;
if pc = 49836 then
	inst <= x"03DC0064";
end if;
if pc = 49840 then
	inst <= x"037E000C";
end if;
if pc = 49844 then
	inst <= x"C57DFFFC";
end if;
if pc = 49848 then
	inst <= x"82003E98";
end if;
if pc = 49852 then
	inst <= x"07DC0064";
end if;
if pc = 49856 then
	inst <= x"C05C0058";
end if;
if pc = 49860 then
	inst <= x"22640220";
end if;
if pc = 49864 then
	inst <= x"C09C0054";
end if;
if pc = 49868 then
	inst <= x"D4286000";
end if;
if pc = 49872 then
	inst <= x"8200C30C";
end if;
if pc = 49876 then
	inst <= x"C51C0054";
end if;
if pc = 49880 then
	inst <= x"C4BC0058";
end if;
if pc = 49884 then
	inst <= x"C17DFFFC";
end if;
if pc = 49888 then
	inst <= x"004E0000";
end if;
if pc = 49892 then
	inst <= x"00320000";
end if;
if pc = 49896 then
	inst <= x"03DC0064";
end if;
if pc = 49900 then
	inst <= x"037E000C";
end if;
if pc = 49904 then
	inst <= x"C57DFFFC";
end if;
if pc = 49908 then
	inst <= x"82003CC4";
end if;
if pc = 49912 then
	inst <= x"07DC0064";
end if;
if pc = 49916 then
	inst <= x"C05C0058";
end if;
if pc = 49920 then
	inst <= x"22640220";
end if;
if pc = 49924 then
	inst <= x"C09C0054";
end if;
if pc = 49928 then
	inst <= x"D4286000";
end if;
if pc = 49932 then
	inst <= x"06240001";
end if;
if pc = 49936 then
	inst <= x"8620C408";
end if;
if pc = 49940 then
	inst <= x"22420220";
end if;
if pc = 49944 then
	inst <= x"C07C0050";
end if;
if pc = 49948 then
	inst <= x"D0464000";
end if;
if pc = 49952 then
	inst <= x"C07C004C";
end if;
if pc = 49956 then
	inst <= x"C0860004";
end if;
if pc = 49960 then
	inst <= x"C0A60000";
end if;
if pc = 49964 then
	inst <= x"C0C40004";
end if;
if pc = 49968 then
	inst <= x"02E00001";
end if;
if pc = 49972 then
	inst <= x"82CEC3B0";
end if;
if pc = 49976 then
	inst <= x"02E00002";
end if;
if pc = 49980 then
	inst <= x"82CEC378";
end if;
if pc = 49984 then
	inst <= x"C49C005C";
end if;
if pc = 49988 then
	inst <= x"C43C0060";
end if;
if pc = 49992 then
	inst <= x"C17DFFFC";
end if;
if pc = 49996 then
	inst <= x"002A0000";
end if;
if pc = 50000 then
	inst <= x"03DC006C";
end if;
if pc = 50004 then
	inst <= x"037E000C";
end if;
if pc = 50008 then
	inst <= x"C57DFFFC";
end if;
if pc = 50012 then
	inst <= x"8200400C";
end if;
if pc = 50016 then
	inst <= x"07DC006C";
end if;
if pc = 50020 then
	inst <= x"C05C0060";
end if;
if pc = 50024 then
	inst <= x"22640220";
end if;
if pc = 50028 then
	inst <= x"C09C005C";
end if;
if pc = 50032 then
	inst <= x"D4286000";
end if;
if pc = 50036 then
	inst <= x"8200C3AC";
end if;
if pc = 50040 then
	inst <= x"C49C005C";
end if;
if pc = 50044 then
	inst <= x"C43C0060";
end if;
if pc = 50048 then
	inst <= x"C17DFFFC";
end if;
if pc = 50052 then
	inst <= x"002A0000";
end if;
if pc = 50056 then
	inst <= x"03DC006C";
end if;
if pc = 50060 then
	inst <= x"037E000C";
end if;
if pc = 50064 then
	inst <= x"C57DFFFC";
end if;
if pc = 50068 then
	inst <= x"82003E98";
end if;
if pc = 50072 then
	inst <= x"07DC006C";
end if;
if pc = 50076 then
	inst <= x"C05C0060";
end if;
if pc = 50080 then
	inst <= x"22640220";
end if;
if pc = 50084 then
	inst <= x"C09C005C";
end if;
if pc = 50088 then
	inst <= x"D4286000";
end if;
if pc = 50092 then
	inst <= x"8200C3E4";
end if;
if pc = 50096 then
	inst <= x"C49C005C";
end if;
if pc = 50100 then
	inst <= x"C43C0060";
end if;
if pc = 50104 then
	inst <= x"C17DFFFC";
end if;
if pc = 50108 then
	inst <= x"002A0000";
end if;
if pc = 50112 then
	inst <= x"03DC006C";
end if;
if pc = 50116 then
	inst <= x"037E000C";
end if;
if pc = 50120 then
	inst <= x"C57DFFFC";
end if;
if pc = 50124 then
	inst <= x"82003CC4";
end if;
if pc = 50128 then
	inst <= x"07DC006C";
end if;
if pc = 50132 then
	inst <= x"C05C0060";
end if;
if pc = 50136 then
	inst <= x"22640220";
end if;
if pc = 50140 then
	inst <= x"C09C005C";
end if;
if pc = 50144 then
	inst <= x"D4286000";
end if;
if pc = 50148 then
	inst <= x"06440001";
end if;
if pc = 50152 then
	inst <= x"C03C004C";
end if;
if pc = 50156 then
	inst <= x"C17DFFFC";
end if;
if pc = 50160 then
	inst <= x"03DC006C";
end if;
if pc = 50164 then
	inst <= x"037E000C";
end if;
if pc = 50168 then
	inst <= x"C57DFFFC";
end if;
if pc = 50172 then
	inst <= x"820042A4";
end if;
if pc = 50176 then
	inst <= x"07DC006C";
end if;
if pc = 50180 then
	inst <= x"8200C408";
end if;
if pc = 50184 then
	inst <= x"8200C40C";
end if;
if pc = 50188 then
	inst <= x"C03C0048";
end if;
if pc = 50192 then
	inst <= x"06220001";
end if;
if pc = 50196 then
	inst <= x"8620C704";
end if;
if pc = 50200 then
	inst <= x"22420220";
end if;
if pc = 50204 then
	inst <= x"C07C0004";
end if;
if pc = 50208 then
	inst <= x"D0464000";
end if;
if pc = 50212 then
	inst <= x"C09C0000";
end if;
if pc = 50216 then
	inst <= x"C0880000";
end if;
if pc = 50220 then
	inst <= x"06880001";
end if;
if pc = 50224 then
	inst <= x"C43C0064";
end if;
if pc = 50228 then
	inst <= x"8680C6F4";
end if;
if pc = 50232 then
	inst <= x"02A000C8";
end if;
if pc = 50236 then
	inst <= x"22C80220";
end if;
if pc = 50240 then
	inst <= x"D0CAC000";
end if;
if pc = 50244 then
	inst <= x"C0E40004";
end if;
if pc = 50248 then
	inst <= x"C1040000";
end if;
if pc = 50252 then
	inst <= x"C12C0004";
end if;
if pc = 50256 then
	inst <= x"03400001";
end if;
if pc = 50260 then
	inst <= x"C45C0068";
end if;
if pc = 50264 then
	inst <= x"C4BC006C";
end if;
if pc = 50268 then
	inst <= x"8334C4E0";
end if;
if pc = 50272 then
	inst <= x"03400002";
end if;
if pc = 50276 then
	inst <= x"8334C4A4";
end if;
if pc = 50280 then
	inst <= x"C4FC0070";
end if;
if pc = 50284 then
	inst <= x"C49C0074";
end if;
if pc = 50288 then
	inst <= x"C17DFFFC";
end if;
if pc = 50292 then
	inst <= x"004C0000";
end if;
if pc = 50296 then
	inst <= x"00300000";
end if;
if pc = 50300 then
	inst <= x"03DC0080";
end if;
if pc = 50304 then
	inst <= x"037E000C";
end if;
if pc = 50308 then
	inst <= x"C57DFFFC";
end if;
if pc = 50312 then
	inst <= x"8200400C";
end if;
if pc = 50316 then
	inst <= x"07DC0080";
end if;
if pc = 50320 then
	inst <= x"C05C0074";
end if;
if pc = 50324 then
	inst <= x"22640220";
end if;
if pc = 50328 then
	inst <= x"C09C0070";
end if;
if pc = 50332 then
	inst <= x"D4286000";
end if;
if pc = 50336 then
	inst <= x"8200C4DC";
end if;
if pc = 50340 then
	inst <= x"C4FC0070";
end if;
if pc = 50344 then
	inst <= x"C49C0074";
end if;
if pc = 50348 then
	inst <= x"C17DFFFC";
end if;
if pc = 50352 then
	inst <= x"004C0000";
end if;
if pc = 50356 then
	inst <= x"00300000";
end if;
if pc = 50360 then
	inst <= x"03DC0080";
end if;
if pc = 50364 then
	inst <= x"037E000C";
end if;
if pc = 50368 then
	inst <= x"C57DFFFC";
end if;
if pc = 50372 then
	inst <= x"82003E98";
end if;
if pc = 50376 then
	inst <= x"07DC0080";
end if;
if pc = 50380 then
	inst <= x"C05C0074";
end if;
if pc = 50384 then
	inst <= x"22640220";
end if;
if pc = 50388 then
	inst <= x"C09C0070";
end if;
if pc = 50392 then
	inst <= x"D4286000";
end if;
if pc = 50396 then
	inst <= x"8200C518";
end if;
if pc = 50400 then
	inst <= x"C4FC0070";
end if;
if pc = 50404 then
	inst <= x"C49C0074";
end if;
if pc = 50408 then
	inst <= x"C17DFFFC";
end if;
if pc = 50412 then
	inst <= x"004C0000";
end if;
if pc = 50416 then
	inst <= x"00300000";
end if;
if pc = 50420 then
	inst <= x"03DC0080";
end if;
if pc = 50424 then
	inst <= x"037E000C";
end if;
if pc = 50428 then
	inst <= x"C57DFFFC";
end if;
if pc = 50432 then
	inst <= x"82003CC4";
end if;
if pc = 50436 then
	inst <= x"07DC0080";
end if;
if pc = 50440 then
	inst <= x"C05C0074";
end if;
if pc = 50444 then
	inst <= x"22640220";
end if;
if pc = 50448 then
	inst <= x"C09C0070";
end if;
if pc = 50452 then
	inst <= x"D4286000";
end if;
if pc = 50456 then
	inst <= x"06240001";
end if;
if pc = 50460 then
	inst <= x"8620C6F0";
end if;
if pc = 50464 then
	inst <= x"22420220";
end if;
if pc = 50468 then
	inst <= x"C07C006C";
end if;
if pc = 50472 then
	inst <= x"D0464000";
end if;
if pc = 50476 then
	inst <= x"C09C0068";
end if;
if pc = 50480 then
	inst <= x"C0A80004";
end if;
if pc = 50484 then
	inst <= x"C0C80000";
end if;
if pc = 50488 then
	inst <= x"C0E40004";
end if;
if pc = 50492 then
	inst <= x"03000001";
end if;
if pc = 50496 then
	inst <= x"82F0C5BC";
end if;
if pc = 50500 then
	inst <= x"03000002";
end if;
if pc = 50504 then
	inst <= x"82F0C584";
end if;
if pc = 50508 then
	inst <= x"C4BC0078";
end if;
if pc = 50512 then
	inst <= x"C43C007C";
end if;
if pc = 50516 then
	inst <= x"C17DFFFC";
end if;
if pc = 50520 then
	inst <= x"002C0000";
end if;
if pc = 50524 then
	inst <= x"03DC0088";
end if;
if pc = 50528 then
	inst <= x"037E000C";
end if;
if pc = 50532 then
	inst <= x"C57DFFFC";
end if;
if pc = 50536 then
	inst <= x"8200400C";
end if;
if pc = 50540 then
	inst <= x"07DC0088";
end if;
if pc = 50544 then
	inst <= x"C05C007C";
end if;
if pc = 50548 then
	inst <= x"22640220";
end if;
if pc = 50552 then
	inst <= x"C09C0078";
end if;
if pc = 50556 then
	inst <= x"D4286000";
end if;
if pc = 50560 then
	inst <= x"8200C5B8";
end if;
if pc = 50564 then
	inst <= x"C4BC0078";
end if;
if pc = 50568 then
	inst <= x"C43C007C";
end if;
if pc = 50572 then
	inst <= x"C17DFFFC";
end if;
if pc = 50576 then
	inst <= x"002C0000";
end if;
if pc = 50580 then
	inst <= x"03DC0088";
end if;
if pc = 50584 then
	inst <= x"037E000C";
end if;
if pc = 50588 then
	inst <= x"C57DFFFC";
end if;
if pc = 50592 then
	inst <= x"82003E98";
end if;
if pc = 50596 then
	inst <= x"07DC0088";
end if;
if pc = 50600 then
	inst <= x"C05C007C";
end if;
if pc = 50604 then
	inst <= x"22640220";
end if;
if pc = 50608 then
	inst <= x"C09C0078";
end if;
if pc = 50612 then
	inst <= x"D4286000";
end if;
if pc = 50616 then
	inst <= x"8200C5F0";
end if;
if pc = 50620 then
	inst <= x"C4BC0078";
end if;
if pc = 50624 then
	inst <= x"C43C007C";
end if;
if pc = 50628 then
	inst <= x"C17DFFFC";
end if;
if pc = 50632 then
	inst <= x"002C0000";
end if;
if pc = 50636 then
	inst <= x"03DC0088";
end if;
if pc = 50640 then
	inst <= x"037E000C";
end if;
if pc = 50644 then
	inst <= x"C57DFFFC";
end if;
if pc = 50648 then
	inst <= x"82003CC4";
end if;
if pc = 50652 then
	inst <= x"07DC0088";
end if;
if pc = 50656 then
	inst <= x"C05C007C";
end if;
if pc = 50660 then
	inst <= x"22640220";
end if;
if pc = 50664 then
	inst <= x"C09C0078";
end if;
if pc = 50668 then
	inst <= x"D4286000";
end if;
if pc = 50672 then
	inst <= x"06240001";
end if;
if pc = 50676 then
	inst <= x"8620C6EC";
end if;
if pc = 50680 then
	inst <= x"22420220";
end if;
if pc = 50684 then
	inst <= x"C07C006C";
end if;
if pc = 50688 then
	inst <= x"D0464000";
end if;
if pc = 50692 then
	inst <= x"C07C0068";
end if;
if pc = 50696 then
	inst <= x"C0860004";
end if;
if pc = 50700 then
	inst <= x"C0A60000";
end if;
if pc = 50704 then
	inst <= x"C0C40004";
end if;
if pc = 50708 then
	inst <= x"02E00001";
end if;
if pc = 50712 then
	inst <= x"82CEC694";
end if;
if pc = 50716 then
	inst <= x"02E00002";
end if;
if pc = 50720 then
	inst <= x"82CEC65C";
end if;
if pc = 50724 then
	inst <= x"C49C0080";
end if;
if pc = 50728 then
	inst <= x"C43C0084";
end if;
if pc = 50732 then
	inst <= x"C17DFFFC";
end if;
if pc = 50736 then
	inst <= x"002A0000";
end if;
if pc = 50740 then
	inst <= x"03DC0090";
end if;
if pc = 50744 then
	inst <= x"037E000C";
end if;
if pc = 50748 then
	inst <= x"C57DFFFC";
end if;
if pc = 50752 then
	inst <= x"8200400C";
end if;
if pc = 50756 then
	inst <= x"07DC0090";
end if;
if pc = 50760 then
	inst <= x"C05C0084";
end if;
if pc = 50764 then
	inst <= x"22640220";
end if;
if pc = 50768 then
	inst <= x"C09C0080";
end if;
if pc = 50772 then
	inst <= x"D4286000";
end if;
if pc = 50776 then
	inst <= x"8200C690";
end if;
if pc = 50780 then
	inst <= x"C49C0080";
end if;
if pc = 50784 then
	inst <= x"C43C0084";
end if;
if pc = 50788 then
	inst <= x"C17DFFFC";
end if;
if pc = 50792 then
	inst <= x"002A0000";
end if;
if pc = 50796 then
	inst <= x"03DC0090";
end if;
if pc = 50800 then
	inst <= x"037E000C";
end if;
if pc = 50804 then
	inst <= x"C57DFFFC";
end if;
if pc = 50808 then
	inst <= x"82003E98";
end if;
if pc = 50812 then
	inst <= x"07DC0090";
end if;
if pc = 50816 then
	inst <= x"C05C0084";
end if;
if pc = 50820 then
	inst <= x"22640220";
end if;
if pc = 50824 then
	inst <= x"C09C0080";
end if;
if pc = 50828 then
	inst <= x"D4286000";
end if;
if pc = 50832 then
	inst <= x"8200C6C8";
end if;
if pc = 50836 then
	inst <= x"C49C0080";
end if;
if pc = 50840 then
	inst <= x"C43C0084";
end if;
if pc = 50844 then
	inst <= x"C17DFFFC";
end if;
if pc = 50848 then
	inst <= x"002A0000";
end if;
if pc = 50852 then
	inst <= x"03DC0090";
end if;
if pc = 50856 then
	inst <= x"037E000C";
end if;
if pc = 50860 then
	inst <= x"C57DFFFC";
end if;
if pc = 50864 then
	inst <= x"82003CC4";
end if;
if pc = 50868 then
	inst <= x"07DC0090";
end if;
if pc = 50872 then
	inst <= x"C05C0084";
end if;
if pc = 50876 then
	inst <= x"22640220";
end if;
if pc = 50880 then
	inst <= x"C09C0080";
end if;
if pc = 50884 then
	inst <= x"D4286000";
end if;
if pc = 50888 then
	inst <= x"06440001";
end if;
if pc = 50892 then
	inst <= x"C03C0068";
end if;
if pc = 50896 then
	inst <= x"C17DFFFC";
end if;
if pc = 50900 then
	inst <= x"03DC0090";
end if;
if pc = 50904 then
	inst <= x"037E000C";
end if;
if pc = 50908 then
	inst <= x"C57DFFFC";
end if;
if pc = 50912 then
	inst <= x"820042A4";
end if;
if pc = 50916 then
	inst <= x"07DC0090";
end if;
if pc = 50920 then
	inst <= x"8200C6EC";
end if;
if pc = 50924 then
	inst <= x"8200C6F0";
end if;
if pc = 50928 then
	inst <= x"8200C6F4";
end if;
if pc = 50932 then
	inst <= x"C03C0064";
end if;
if pc = 50936 then
	inst <= x"06420001";
end if;
if pc = 50940 then
	inst <= x"C03C0004";
end if;
if pc = 50944 then
	inst <= x"8200BD10";
end if;
if pc = 50948 then
	inst <= x"C1FDFFFC";
end if;
if pc = 50952 then
	inst <= x"C1FDFFFC";
end if;
if pc = 50956 then
	inst <= x"C1FDFFFC";
end if;
if pc = 50960 then
	inst <= x"C1FDFFFC";
end if;
if pc = 50964 then
	inst <= x"8620D760";
end if;
if pc = 50968 then
	inst <= x"02400354";
end if;
if pc = 50972 then
	inst <= x"22620220";
end if;
if pc = 50976 then
	inst <= x"D0646000";
end if;
if pc = 50980 then
	inst <= x"C08601DC";
end if;
if pc = 50984 then
	inst <= x"02A000C4";
end if;
if pc = 50988 then
	inst <= x"C0CA0000";
end if;
if pc = 50992 then
	inst <= x"06CC0001";
end if;
if pc = 50996 then
	inst <= x"C45C0000";
end if;
if pc = 51000 then
	inst <= x"C43C0004";
end if;
if pc = 51004 then
	inst <= x"C4BC0008";
end if;
if pc = 51008 then
	inst <= x"C47C000C";
end if;
if pc = 51012 then
	inst <= x"86C0CA04";
end if;
if pc = 51016 then
	inst <= x"02E000C8";
end if;
if pc = 51020 then
	inst <= x"230C0220";
end if;
if pc = 51024 then
	inst <= x"D10F0000";
end if;
if pc = 51028 then
	inst <= x"C1280004";
end if;
if pc = 51032 then
	inst <= x"C1480000";
end if;
if pc = 51036 then
	inst <= x"C0500004";
end if;
if pc = 51040 then
	inst <= x"02200001";
end if;
if pc = 51044 then
	inst <= x"C49C0010";
end if;
if pc = 51048 then
	inst <= x"C4FC0014";
end if;
if pc = 51052 then
	inst <= x"8242C7F0";
end if;
if pc = 51056 then
	inst <= x"02200002";
end if;
if pc = 51060 then
	inst <= x"8242C7B4";
end if;
if pc = 51064 then
	inst <= x"C53C0018";
end if;
if pc = 51068 then
	inst <= x"C4DC001C";
end if;
if pc = 51072 then
	inst <= x"C17DFFFC";
end if;
if pc = 51076 then
	inst <= x"00500000";
end if;
if pc = 51080 then
	inst <= x"00340000";
end if;
if pc = 51084 then
	inst <= x"03DC0028";
end if;
if pc = 51088 then
	inst <= x"037E000C";
end if;
if pc = 51092 then
	inst <= x"C57DFFFC";
end if;
if pc = 51096 then
	inst <= x"8200400C";
end if;
if pc = 51100 then
	inst <= x"07DC0028";
end if;
if pc = 51104 then
	inst <= x"C05C001C";
end if;
if pc = 51108 then
	inst <= x"22640220";
end if;
if pc = 51112 then
	inst <= x"C09C0018";
end if;
if pc = 51116 then
	inst <= x"D4286000";
end if;
if pc = 51120 then
	inst <= x"8200C7EC";
end if;
if pc = 51124 then
	inst <= x"C53C0018";
end if;
if pc = 51128 then
	inst <= x"C4DC001C";
end if;
if pc = 51132 then
	inst <= x"C17DFFFC";
end if;
if pc = 51136 then
	inst <= x"00500000";
end if;
if pc = 51140 then
	inst <= x"00340000";
end if;
if pc = 51144 then
	inst <= x"03DC0028";
end if;
if pc = 51148 then
	inst <= x"037E000C";
end if;
if pc = 51152 then
	inst <= x"C57DFFFC";
end if;
if pc = 51156 then
	inst <= x"82003E98";
end if;
if pc = 51160 then
	inst <= x"07DC0028";
end if;
if pc = 51164 then
	inst <= x"C05C001C";
end if;
if pc = 51168 then
	inst <= x"22640220";
end if;
if pc = 51172 then
	inst <= x"C09C0018";
end if;
if pc = 51176 then
	inst <= x"D4286000";
end if;
if pc = 51180 then
	inst <= x"8200C828";
end if;
if pc = 51184 then
	inst <= x"C53C0018";
end if;
if pc = 51188 then
	inst <= x"C4DC001C";
end if;
if pc = 51192 then
	inst <= x"C17DFFFC";
end if;
if pc = 51196 then
	inst <= x"00500000";
end if;
if pc = 51200 then
	inst <= x"00340000";
end if;
if pc = 51204 then
	inst <= x"03DC0028";
end if;
if pc = 51208 then
	inst <= x"037E000C";
end if;
if pc = 51212 then
	inst <= x"C57DFFFC";
end if;
if pc = 51216 then
	inst <= x"82003CC4";
end if;
if pc = 51220 then
	inst <= x"07DC0028";
end if;
if pc = 51224 then
	inst <= x"C05C001C";
end if;
if pc = 51228 then
	inst <= x"22640220";
end if;
if pc = 51232 then
	inst <= x"C09C0018";
end if;
if pc = 51236 then
	inst <= x"D4286000";
end if;
if pc = 51240 then
	inst <= x"06240001";
end if;
if pc = 51244 then
	inst <= x"8620CA00";
end if;
if pc = 51248 then
	inst <= x"22420220";
end if;
if pc = 51252 then
	inst <= x"C07C0014";
end if;
if pc = 51256 then
	inst <= x"D0464000";
end if;
if pc = 51260 then
	inst <= x"C09C0010";
end if;
if pc = 51264 then
	inst <= x"C0A80004";
end if;
if pc = 51268 then
	inst <= x"C0C80000";
end if;
if pc = 51272 then
	inst <= x"C0E40004";
end if;
if pc = 51276 then
	inst <= x"03000001";
end if;
if pc = 51280 then
	inst <= x"82F0C8CC";
end if;
if pc = 51284 then
	inst <= x"03000002";
end if;
if pc = 51288 then
	inst <= x"82F0C894";
end if;
if pc = 51292 then
	inst <= x"C4BC0020";
end if;
if pc = 51296 then
	inst <= x"C43C0024";
end if;
if pc = 51300 then
	inst <= x"C17DFFFC";
end if;
if pc = 51304 then
	inst <= x"002C0000";
end if;
if pc = 51308 then
	inst <= x"03DC0030";
end if;
if pc = 51312 then
	inst <= x"037E000C";
end if;
if pc = 51316 then
	inst <= x"C57DFFFC";
end if;
if pc = 51320 then
	inst <= x"8200400C";
end if;
if pc = 51324 then
	inst <= x"07DC0030";
end if;
if pc = 51328 then
	inst <= x"C05C0024";
end if;
if pc = 51332 then
	inst <= x"22640220";
end if;
if pc = 51336 then
	inst <= x"C09C0020";
end if;
if pc = 51340 then
	inst <= x"D4286000";
end if;
if pc = 51344 then
	inst <= x"8200C8C8";
end if;
if pc = 51348 then
	inst <= x"C4BC0020";
end if;
if pc = 51352 then
	inst <= x"C43C0024";
end if;
if pc = 51356 then
	inst <= x"C17DFFFC";
end if;
if pc = 51360 then
	inst <= x"002C0000";
end if;
if pc = 51364 then
	inst <= x"03DC0030";
end if;
if pc = 51368 then
	inst <= x"037E000C";
end if;
if pc = 51372 then
	inst <= x"C57DFFFC";
end if;
if pc = 51376 then
	inst <= x"82003E98";
end if;
if pc = 51380 then
	inst <= x"07DC0030";
end if;
if pc = 51384 then
	inst <= x"C05C0024";
end if;
if pc = 51388 then
	inst <= x"22640220";
end if;
if pc = 51392 then
	inst <= x"C09C0020";
end if;
if pc = 51396 then
	inst <= x"D4286000";
end if;
if pc = 51400 then
	inst <= x"8200C900";
end if;
if pc = 51404 then
	inst <= x"C4BC0020";
end if;
if pc = 51408 then
	inst <= x"C43C0024";
end if;
if pc = 51412 then
	inst <= x"C17DFFFC";
end if;
if pc = 51416 then
	inst <= x"002C0000";
end if;
if pc = 51420 then
	inst <= x"03DC0030";
end if;
if pc = 51424 then
	inst <= x"037E000C";
end if;
if pc = 51428 then
	inst <= x"C57DFFFC";
end if;
if pc = 51432 then
	inst <= x"82003CC4";
end if;
if pc = 51436 then
	inst <= x"07DC0030";
end if;
if pc = 51440 then
	inst <= x"C05C0024";
end if;
if pc = 51444 then
	inst <= x"22640220";
end if;
if pc = 51448 then
	inst <= x"C09C0020";
end if;
if pc = 51452 then
	inst <= x"D4286000";
end if;
if pc = 51456 then
	inst <= x"06240001";
end if;
if pc = 51460 then
	inst <= x"8620C9FC";
end if;
if pc = 51464 then
	inst <= x"22420220";
end if;
if pc = 51468 then
	inst <= x"C07C0014";
end if;
if pc = 51472 then
	inst <= x"D0464000";
end if;
if pc = 51476 then
	inst <= x"C07C0010";
end if;
if pc = 51480 then
	inst <= x"C0860004";
end if;
if pc = 51484 then
	inst <= x"C0A60000";
end if;
if pc = 51488 then
	inst <= x"C0C40004";
end if;
if pc = 51492 then
	inst <= x"02E00001";
end if;
if pc = 51496 then
	inst <= x"82CEC9A4";
end if;
if pc = 51500 then
	inst <= x"02E00002";
end if;
if pc = 51504 then
	inst <= x"82CEC96C";
end if;
if pc = 51508 then
	inst <= x"C49C0028";
end if;
if pc = 51512 then
	inst <= x"C43C002C";
end if;
if pc = 51516 then
	inst <= x"C17DFFFC";
end if;
if pc = 51520 then
	inst <= x"002A0000";
end if;
if pc = 51524 then
	inst <= x"03DC0038";
end if;
if pc = 51528 then
	inst <= x"037E000C";
end if;
if pc = 51532 then
	inst <= x"C57DFFFC";
end if;
if pc = 51536 then
	inst <= x"8200400C";
end if;
if pc = 51540 then
	inst <= x"07DC0038";
end if;
if pc = 51544 then
	inst <= x"C05C002C";
end if;
if pc = 51548 then
	inst <= x"22640220";
end if;
if pc = 51552 then
	inst <= x"C09C0028";
end if;
if pc = 51556 then
	inst <= x"D4286000";
end if;
if pc = 51560 then
	inst <= x"8200C9A0";
end if;
if pc = 51564 then
	inst <= x"C49C0028";
end if;
if pc = 51568 then
	inst <= x"C43C002C";
end if;
if pc = 51572 then
	inst <= x"C17DFFFC";
end if;
if pc = 51576 then
	inst <= x"002A0000";
end if;
if pc = 51580 then
	inst <= x"03DC0038";
end if;
if pc = 51584 then
	inst <= x"037E000C";
end if;
if pc = 51588 then
	inst <= x"C57DFFFC";
end if;
if pc = 51592 then
	inst <= x"82003E98";
end if;
if pc = 51596 then
	inst <= x"07DC0038";
end if;
if pc = 51600 then
	inst <= x"C05C002C";
end if;
if pc = 51604 then
	inst <= x"22640220";
end if;
if pc = 51608 then
	inst <= x"C09C0028";
end if;
if pc = 51612 then
	inst <= x"D4286000";
end if;
if pc = 51616 then
	inst <= x"8200C9D8";
end if;
if pc = 51620 then
	inst <= x"C49C0028";
end if;
if pc = 51624 then
	inst <= x"C43C002C";
end if;
if pc = 51628 then
	inst <= x"C17DFFFC";
end if;
if pc = 51632 then
	inst <= x"002A0000";
end if;
if pc = 51636 then
	inst <= x"03DC0038";
end if;
if pc = 51640 then
	inst <= x"037E000C";
end if;
if pc = 51644 then
	inst <= x"C57DFFFC";
end if;
if pc = 51648 then
	inst <= x"82003CC4";
end if;
if pc = 51652 then
	inst <= x"07DC0038";
end if;
if pc = 51656 then
	inst <= x"C05C002C";
end if;
if pc = 51660 then
	inst <= x"22640220";
end if;
if pc = 51664 then
	inst <= x"C09C0028";
end if;
if pc = 51668 then
	inst <= x"D4286000";
end if;
if pc = 51672 then
	inst <= x"06440001";
end if;
if pc = 51676 then
	inst <= x"C03C0010";
end if;
if pc = 51680 then
	inst <= x"C17DFFFC";
end if;
if pc = 51684 then
	inst <= x"03DC0038";
end if;
if pc = 51688 then
	inst <= x"037E000C";
end if;
if pc = 51692 then
	inst <= x"C57DFFFC";
end if;
if pc = 51696 then
	inst <= x"820042A4";
end if;
if pc = 51700 then
	inst <= x"07DC0038";
end if;
if pc = 51704 then
	inst <= x"8200C9FC";
end if;
if pc = 51708 then
	inst <= x"8200CA00";
end if;
if pc = 51712 then
	inst <= x"8200CA04";
end if;
if pc = 51716 then
	inst <= x"C03C000C";
end if;
if pc = 51720 then
	inst <= x"C04201D8";
end if;
if pc = 51724 then
	inst <= x"C07C0008";
end if;
if pc = 51728 then
	inst <= x"C0860000";
end if;
if pc = 51732 then
	inst <= x"06880001";
end if;
if pc = 51736 then
	inst <= x"8680CBFC";
end if;
if pc = 51740 then
	inst <= x"02A000C8";
end if;
if pc = 51744 then
	inst <= x"22C80220";
end if;
if pc = 51748 then
	inst <= x"D0CAC000";
end if;
if pc = 51752 then
	inst <= x"C0E40004";
end if;
if pc = 51756 then
	inst <= x"C1040000";
end if;
if pc = 51760 then
	inst <= x"C12C0004";
end if;
if pc = 51764 then
	inst <= x"03400001";
end if;
if pc = 51768 then
	inst <= x"C45C0030";
end if;
if pc = 51772 then
	inst <= x"C4BC0034";
end if;
if pc = 51776 then
	inst <= x"8334CAC4";
end if;
if pc = 51780 then
	inst <= x"03400002";
end if;
if pc = 51784 then
	inst <= x"8334CA88";
end if;
if pc = 51788 then
	inst <= x"C4FC0038";
end if;
if pc = 51792 then
	inst <= x"C49C003C";
end if;
if pc = 51796 then
	inst <= x"C17DFFFC";
end if;
if pc = 51800 then
	inst <= x"004C0000";
end if;
if pc = 51804 then
	inst <= x"00300000";
end if;
if pc = 51808 then
	inst <= x"03DC0048";
end if;
if pc = 51812 then
	inst <= x"037E000C";
end if;
if pc = 51816 then
	inst <= x"C57DFFFC";
end if;
if pc = 51820 then
	inst <= x"8200400C";
end if;
if pc = 51824 then
	inst <= x"07DC0048";
end if;
if pc = 51828 then
	inst <= x"C05C003C";
end if;
if pc = 51832 then
	inst <= x"22640220";
end if;
if pc = 51836 then
	inst <= x"C09C0038";
end if;
if pc = 51840 then
	inst <= x"D4286000";
end if;
if pc = 51844 then
	inst <= x"8200CAC0";
end if;
if pc = 51848 then
	inst <= x"C4FC0038";
end if;
if pc = 51852 then
	inst <= x"C49C003C";
end if;
if pc = 51856 then
	inst <= x"C17DFFFC";
end if;
if pc = 51860 then
	inst <= x"004C0000";
end if;
if pc = 51864 then
	inst <= x"00300000";
end if;
if pc = 51868 then
	inst <= x"03DC0048";
end if;
if pc = 51872 then
	inst <= x"037E000C";
end if;
if pc = 51876 then
	inst <= x"C57DFFFC";
end if;
if pc = 51880 then
	inst <= x"82003E98";
end if;
if pc = 51884 then
	inst <= x"07DC0048";
end if;
if pc = 51888 then
	inst <= x"C05C003C";
end if;
if pc = 51892 then
	inst <= x"22640220";
end if;
if pc = 51896 then
	inst <= x"C09C0038";
end if;
if pc = 51900 then
	inst <= x"D4286000";
end if;
if pc = 51904 then
	inst <= x"8200CAFC";
end if;
if pc = 51908 then
	inst <= x"C4FC0038";
end if;
if pc = 51912 then
	inst <= x"C49C003C";
end if;
if pc = 51916 then
	inst <= x"C17DFFFC";
end if;
if pc = 51920 then
	inst <= x"004C0000";
end if;
if pc = 51924 then
	inst <= x"00300000";
end if;
if pc = 51928 then
	inst <= x"03DC0048";
end if;
if pc = 51932 then
	inst <= x"037E000C";
end if;
if pc = 51936 then
	inst <= x"C57DFFFC";
end if;
if pc = 51940 then
	inst <= x"82003CC4";
end if;
if pc = 51944 then
	inst <= x"07DC0048";
end if;
if pc = 51948 then
	inst <= x"C05C003C";
end if;
if pc = 51952 then
	inst <= x"22640220";
end if;
if pc = 51956 then
	inst <= x"C09C0038";
end if;
if pc = 51960 then
	inst <= x"D4286000";
end if;
if pc = 51964 then
	inst <= x"06240001";
end if;
if pc = 51968 then
	inst <= x"8620CBF8";
end if;
if pc = 51972 then
	inst <= x"22420220";
end if;
if pc = 51976 then
	inst <= x"C07C0034";
end if;
if pc = 51980 then
	inst <= x"D0464000";
end if;
if pc = 51984 then
	inst <= x"C07C0030";
end if;
if pc = 51988 then
	inst <= x"C0860004";
end if;
if pc = 51992 then
	inst <= x"C0A60000";
end if;
if pc = 51996 then
	inst <= x"C0C40004";
end if;
if pc = 52000 then
	inst <= x"02E00001";
end if;
if pc = 52004 then
	inst <= x"82CECBA0";
end if;
if pc = 52008 then
	inst <= x"02E00002";
end if;
if pc = 52012 then
	inst <= x"82CECB68";
end if;
if pc = 52016 then
	inst <= x"C49C0040";
end if;
if pc = 52020 then
	inst <= x"C43C0044";
end if;
if pc = 52024 then
	inst <= x"C17DFFFC";
end if;
if pc = 52028 then
	inst <= x"002A0000";
end if;
if pc = 52032 then
	inst <= x"03DC0050";
end if;
if pc = 52036 then
	inst <= x"037E000C";
end if;
if pc = 52040 then
	inst <= x"C57DFFFC";
end if;
if pc = 52044 then
	inst <= x"8200400C";
end if;
if pc = 52048 then
	inst <= x"07DC0050";
end if;
if pc = 52052 then
	inst <= x"C05C0044";
end if;
if pc = 52056 then
	inst <= x"22640220";
end if;
if pc = 52060 then
	inst <= x"C09C0040";
end if;
if pc = 52064 then
	inst <= x"D4286000";
end if;
if pc = 52068 then
	inst <= x"8200CB9C";
end if;
if pc = 52072 then
	inst <= x"C49C0040";
end if;
if pc = 52076 then
	inst <= x"C43C0044";
end if;
if pc = 52080 then
	inst <= x"C17DFFFC";
end if;
if pc = 52084 then
	inst <= x"002A0000";
end if;
if pc = 52088 then
	inst <= x"03DC0050";
end if;
if pc = 52092 then
	inst <= x"037E000C";
end if;
if pc = 52096 then
	inst <= x"C57DFFFC";
end if;
if pc = 52100 then
	inst <= x"82003E98";
end if;
if pc = 52104 then
	inst <= x"07DC0050";
end if;
if pc = 52108 then
	inst <= x"C05C0044";
end if;
if pc = 52112 then
	inst <= x"22640220";
end if;
if pc = 52116 then
	inst <= x"C09C0040";
end if;
if pc = 52120 then
	inst <= x"D4286000";
end if;
if pc = 52124 then
	inst <= x"8200CBD4";
end if;
if pc = 52128 then
	inst <= x"C49C0040";
end if;
if pc = 52132 then
	inst <= x"C43C0044";
end if;
if pc = 52136 then
	inst <= x"C17DFFFC";
end if;
if pc = 52140 then
	inst <= x"002A0000";
end if;
if pc = 52144 then
	inst <= x"03DC0050";
end if;
if pc = 52148 then
	inst <= x"037E000C";
end if;
if pc = 52152 then
	inst <= x"C57DFFFC";
end if;
if pc = 52156 then
	inst <= x"82003CC4";
end if;
if pc = 52160 then
	inst <= x"07DC0050";
end if;
if pc = 52164 then
	inst <= x"C05C0044";
end if;
if pc = 52168 then
	inst <= x"22640220";
end if;
if pc = 52172 then
	inst <= x"C09C0040";
end if;
if pc = 52176 then
	inst <= x"D4286000";
end if;
if pc = 52180 then
	inst <= x"06440001";
end if;
if pc = 52184 then
	inst <= x"C03C0030";
end if;
if pc = 52188 then
	inst <= x"C17DFFFC";
end if;
if pc = 52192 then
	inst <= x"03DC0050";
end if;
if pc = 52196 then
	inst <= x"037E000C";
end if;
if pc = 52200 then
	inst <= x"C57DFFFC";
end if;
if pc = 52204 then
	inst <= x"820042A4";
end if;
if pc = 52208 then
	inst <= x"07DC0050";
end if;
if pc = 52212 then
	inst <= x"8200CBF8";
end if;
if pc = 52216 then
	inst <= x"8200CBFC";
end if;
if pc = 52220 then
	inst <= x"C03C000C";
end if;
if pc = 52224 then
	inst <= x"C04201D4";
end if;
if pc = 52228 then
	inst <= x"C07C0008";
end if;
if pc = 52232 then
	inst <= x"C0860000";
end if;
if pc = 52236 then
	inst <= x"06880001";
end if;
if pc = 52240 then
	inst <= x"8680CED0";
end if;
if pc = 52244 then
	inst <= x"02A000C8";
end if;
if pc = 52248 then
	inst <= x"22C80220";
end if;
if pc = 52252 then
	inst <= x"D0CAC000";
end if;
if pc = 52256 then
	inst <= x"C0E40004";
end if;
if pc = 52260 then
	inst <= x"C1040000";
end if;
if pc = 52264 then
	inst <= x"C12C0004";
end if;
if pc = 52268 then
	inst <= x"03400001";
end if;
if pc = 52272 then
	inst <= x"C45C0048";
end if;
if pc = 52276 then
	inst <= x"C4BC004C";
end if;
if pc = 52280 then
	inst <= x"8334CCBC";
end if;
if pc = 52284 then
	inst <= x"03400002";
end if;
if pc = 52288 then
	inst <= x"8334CC80";
end if;
if pc = 52292 then
	inst <= x"C4FC0050";
end if;
if pc = 52296 then
	inst <= x"C49C0054";
end if;
if pc = 52300 then
	inst <= x"C17DFFFC";
end if;
if pc = 52304 then
	inst <= x"004C0000";
end if;
if pc = 52308 then
	inst <= x"00300000";
end if;
if pc = 52312 then
	inst <= x"03DC0060";
end if;
if pc = 52316 then
	inst <= x"037E000C";
end if;
if pc = 52320 then
	inst <= x"C57DFFFC";
end if;
if pc = 52324 then
	inst <= x"8200400C";
end if;
if pc = 52328 then
	inst <= x"07DC0060";
end if;
if pc = 52332 then
	inst <= x"C05C0054";
end if;
if pc = 52336 then
	inst <= x"22640220";
end if;
if pc = 52340 then
	inst <= x"C09C0050";
end if;
if pc = 52344 then
	inst <= x"D4286000";
end if;
if pc = 52348 then
	inst <= x"8200CCB8";
end if;
if pc = 52352 then
	inst <= x"C4FC0050";
end if;
if pc = 52356 then
	inst <= x"C49C0054";
end if;
if pc = 52360 then
	inst <= x"C17DFFFC";
end if;
if pc = 52364 then
	inst <= x"004C0000";
end if;
if pc = 52368 then
	inst <= x"00300000";
end if;
if pc = 52372 then
	inst <= x"03DC0060";
end if;
if pc = 52376 then
	inst <= x"037E000C";
end if;
if pc = 52380 then
	inst <= x"C57DFFFC";
end if;
if pc = 52384 then
	inst <= x"82003E98";
end if;
if pc = 52388 then
	inst <= x"07DC0060";
end if;
if pc = 52392 then
	inst <= x"C05C0054";
end if;
if pc = 52396 then
	inst <= x"22640220";
end if;
if pc = 52400 then
	inst <= x"C09C0050";
end if;
if pc = 52404 then
	inst <= x"D4286000";
end if;
if pc = 52408 then
	inst <= x"8200CCF4";
end if;
if pc = 52412 then
	inst <= x"C4FC0050";
end if;
if pc = 52416 then
	inst <= x"C49C0054";
end if;
if pc = 52420 then
	inst <= x"C17DFFFC";
end if;
if pc = 52424 then
	inst <= x"004C0000";
end if;
if pc = 52428 then
	inst <= x"00300000";
end if;
if pc = 52432 then
	inst <= x"03DC0060";
end if;
if pc = 52436 then
	inst <= x"037E000C";
end if;
if pc = 52440 then
	inst <= x"C57DFFFC";
end if;
if pc = 52444 then
	inst <= x"82003CC4";
end if;
if pc = 52448 then
	inst <= x"07DC0060";
end if;
if pc = 52452 then
	inst <= x"C05C0054";
end if;
if pc = 52456 then
	inst <= x"22640220";
end if;
if pc = 52460 then
	inst <= x"C09C0050";
end if;
if pc = 52464 then
	inst <= x"D4286000";
end if;
if pc = 52468 then
	inst <= x"06240001";
end if;
if pc = 52472 then
	inst <= x"8620CECC";
end if;
if pc = 52476 then
	inst <= x"22420220";
end if;
if pc = 52480 then
	inst <= x"C07C004C";
end if;
if pc = 52484 then
	inst <= x"D0464000";
end if;
if pc = 52488 then
	inst <= x"C09C0048";
end if;
if pc = 52492 then
	inst <= x"C0A80004";
end if;
if pc = 52496 then
	inst <= x"C0C80000";
end if;
if pc = 52500 then
	inst <= x"C0E40004";
end if;
if pc = 52504 then
	inst <= x"03000001";
end if;
if pc = 52508 then
	inst <= x"82F0CD98";
end if;
if pc = 52512 then
	inst <= x"03000002";
end if;
if pc = 52516 then
	inst <= x"82F0CD60";
end if;
if pc = 52520 then
	inst <= x"C4BC0058";
end if;
if pc = 52524 then
	inst <= x"C43C005C";
end if;
if pc = 52528 then
	inst <= x"C17DFFFC";
end if;
if pc = 52532 then
	inst <= x"002C0000";
end if;
if pc = 52536 then
	inst <= x"03DC0068";
end if;
if pc = 52540 then
	inst <= x"037E000C";
end if;
if pc = 52544 then
	inst <= x"C57DFFFC";
end if;
if pc = 52548 then
	inst <= x"8200400C";
end if;
if pc = 52552 then
	inst <= x"07DC0068";
end if;
if pc = 52556 then
	inst <= x"C05C005C";
end if;
if pc = 52560 then
	inst <= x"22640220";
end if;
if pc = 52564 then
	inst <= x"C09C0058";
end if;
if pc = 52568 then
	inst <= x"D4286000";
end if;
if pc = 52572 then
	inst <= x"8200CD94";
end if;
if pc = 52576 then
	inst <= x"C4BC0058";
end if;
if pc = 52580 then
	inst <= x"C43C005C";
end if;
if pc = 52584 then
	inst <= x"C17DFFFC";
end if;
if pc = 52588 then
	inst <= x"002C0000";
end if;
if pc = 52592 then
	inst <= x"03DC0068";
end if;
if pc = 52596 then
	inst <= x"037E000C";
end if;
if pc = 52600 then
	inst <= x"C57DFFFC";
end if;
if pc = 52604 then
	inst <= x"82003E98";
end if;
if pc = 52608 then
	inst <= x"07DC0068";
end if;
if pc = 52612 then
	inst <= x"C05C005C";
end if;
if pc = 52616 then
	inst <= x"22640220";
end if;
if pc = 52620 then
	inst <= x"C09C0058";
end if;
if pc = 52624 then
	inst <= x"D4286000";
end if;
if pc = 52628 then
	inst <= x"8200CDCC";
end if;
if pc = 52632 then
	inst <= x"C4BC0058";
end if;
if pc = 52636 then
	inst <= x"C43C005C";
end if;
if pc = 52640 then
	inst <= x"C17DFFFC";
end if;
if pc = 52644 then
	inst <= x"002C0000";
end if;
if pc = 52648 then
	inst <= x"03DC0068";
end if;
if pc = 52652 then
	inst <= x"037E000C";
end if;
if pc = 52656 then
	inst <= x"C57DFFFC";
end if;
if pc = 52660 then
	inst <= x"82003CC4";
end if;
if pc = 52664 then
	inst <= x"07DC0068";
end if;
if pc = 52668 then
	inst <= x"C05C005C";
end if;
if pc = 52672 then
	inst <= x"22640220";
end if;
if pc = 52676 then
	inst <= x"C09C0058";
end if;
if pc = 52680 then
	inst <= x"D4286000";
end if;
if pc = 52684 then
	inst <= x"06240001";
end if;
if pc = 52688 then
	inst <= x"8620CEC8";
end if;
if pc = 52692 then
	inst <= x"22420220";
end if;
if pc = 52696 then
	inst <= x"C07C004C";
end if;
if pc = 52700 then
	inst <= x"D0464000";
end if;
if pc = 52704 then
	inst <= x"C07C0048";
end if;
if pc = 52708 then
	inst <= x"C0860004";
end if;
if pc = 52712 then
	inst <= x"C0A60000";
end if;
if pc = 52716 then
	inst <= x"C0C40004";
end if;
if pc = 52720 then
	inst <= x"02E00001";
end if;
if pc = 52724 then
	inst <= x"82CECE70";
end if;
if pc = 52728 then
	inst <= x"02E00002";
end if;
if pc = 52732 then
	inst <= x"82CECE38";
end if;
if pc = 52736 then
	inst <= x"C49C0060";
end if;
if pc = 52740 then
	inst <= x"C43C0064";
end if;
if pc = 52744 then
	inst <= x"C17DFFFC";
end if;
if pc = 52748 then
	inst <= x"002A0000";
end if;
if pc = 52752 then
	inst <= x"03DC0070";
end if;
if pc = 52756 then
	inst <= x"037E000C";
end if;
if pc = 52760 then
	inst <= x"C57DFFFC";
end if;
if pc = 52764 then
	inst <= x"8200400C";
end if;
if pc = 52768 then
	inst <= x"07DC0070";
end if;
if pc = 52772 then
	inst <= x"C05C0064";
end if;
if pc = 52776 then
	inst <= x"22640220";
end if;
if pc = 52780 then
	inst <= x"C09C0060";
end if;
if pc = 52784 then
	inst <= x"D4286000";
end if;
if pc = 52788 then
	inst <= x"8200CE6C";
end if;
if pc = 52792 then
	inst <= x"C49C0060";
end if;
if pc = 52796 then
	inst <= x"C43C0064";
end if;
if pc = 52800 then
	inst <= x"C17DFFFC";
end if;
if pc = 52804 then
	inst <= x"002A0000";
end if;
if pc = 52808 then
	inst <= x"03DC0070";
end if;
if pc = 52812 then
	inst <= x"037E000C";
end if;
if pc = 52816 then
	inst <= x"C57DFFFC";
end if;
if pc = 52820 then
	inst <= x"82003E98";
end if;
if pc = 52824 then
	inst <= x"07DC0070";
end if;
if pc = 52828 then
	inst <= x"C05C0064";
end if;
if pc = 52832 then
	inst <= x"22640220";
end if;
if pc = 52836 then
	inst <= x"C09C0060";
end if;
if pc = 52840 then
	inst <= x"D4286000";
end if;
if pc = 52844 then
	inst <= x"8200CEA4";
end if;
if pc = 52848 then
	inst <= x"C49C0060";
end if;
if pc = 52852 then
	inst <= x"C43C0064";
end if;
if pc = 52856 then
	inst <= x"C17DFFFC";
end if;
if pc = 52860 then
	inst <= x"002A0000";
end if;
if pc = 52864 then
	inst <= x"03DC0070";
end if;
if pc = 52868 then
	inst <= x"037E000C";
end if;
if pc = 52872 then
	inst <= x"C57DFFFC";
end if;
if pc = 52876 then
	inst <= x"82003CC4";
end if;
if pc = 52880 then
	inst <= x"07DC0070";
end if;
if pc = 52884 then
	inst <= x"C05C0064";
end if;
if pc = 52888 then
	inst <= x"22640220";
end if;
if pc = 52892 then
	inst <= x"C09C0060";
end if;
if pc = 52896 then
	inst <= x"D4286000";
end if;
if pc = 52900 then
	inst <= x"06440001";
end if;
if pc = 52904 then
	inst <= x"C03C0048";
end if;
if pc = 52908 then
	inst <= x"C17DFFFC";
end if;
if pc = 52912 then
	inst <= x"03DC0070";
end if;
if pc = 52916 then
	inst <= x"037E000C";
end if;
if pc = 52920 then
	inst <= x"C57DFFFC";
end if;
if pc = 52924 then
	inst <= x"820042A4";
end if;
if pc = 52928 then
	inst <= x"07DC0070";
end if;
if pc = 52932 then
	inst <= x"8200CEC8";
end if;
if pc = 52936 then
	inst <= x"8200CECC";
end if;
if pc = 52940 then
	inst <= x"8200CED0";
end if;
if pc = 52944 then
	inst <= x"02400074";
end if;
if pc = 52948 then
	inst <= x"C03C000C";
end if;
if pc = 52952 then
	inst <= x"C17DFFFC";
end if;
if pc = 52956 then
	inst <= x"03DC0070";
end if;
if pc = 52960 then
	inst <= x"037E000C";
end if;
if pc = 52964 then
	inst <= x"C57DFFFC";
end if;
if pc = 52968 then
	inst <= x"8200BD10";
end if;
if pc = 52972 then
	inst <= x"07DC0070";
end if;
if pc = 52976 then
	inst <= x"C03C0004";
end if;
if pc = 52980 then
	inst <= x"06220001";
end if;
if pc = 52984 then
	inst <= x"8620D75C";
end if;
if pc = 52988 then
	inst <= x"22420220";
end if;
if pc = 52992 then
	inst <= x"C07C0000";
end if;
if pc = 52996 then
	inst <= x"D0464000";
end if;
if pc = 53000 then
	inst <= x"C08401DC";
end if;
if pc = 53004 then
	inst <= x"C0BC0008";
end if;
if pc = 53008 then
	inst <= x"C0CA0000";
end if;
if pc = 53012 then
	inst <= x"06CC0001";
end if;
if pc = 53016 then
	inst <= x"C43C0068";
end if;
if pc = 53020 then
	inst <= x"C45C006C";
end if;
if pc = 53024 then
	inst <= x"86C0D104";
end if;
if pc = 53028 then
	inst <= x"02E000C8";
end if;
if pc = 53032 then
	inst <= x"230C0220";
end if;
if pc = 53036 then
	inst <= x"D10F0000";
end if;
if pc = 53040 then
	inst <= x"C1280004";
end if;
if pc = 53044 then
	inst <= x"C1480000";
end if;
if pc = 53048 then
	inst <= x"C0700004";
end if;
if pc = 53052 then
	inst <= x"02200001";
end if;
if pc = 53056 then
	inst <= x"C49C0070";
end if;
if pc = 53060 then
	inst <= x"C4FC0074";
end if;
if pc = 53064 then
	inst <= x"8262CFCC";
end if;
if pc = 53068 then
	inst <= x"02200002";
end if;
if pc = 53072 then
	inst <= x"8262CF90";
end if;
if pc = 53076 then
	inst <= x"C53C0078";
end if;
if pc = 53080 then
	inst <= x"C4DC007C";
end if;
if pc = 53084 then
	inst <= x"C17DFFFC";
end if;
if pc = 53088 then
	inst <= x"00500000";
end if;
if pc = 53092 then
	inst <= x"00340000";
end if;
if pc = 53096 then
	inst <= x"03DC0088";
end if;
if pc = 53100 then
	inst <= x"037E000C";
end if;
if pc = 53104 then
	inst <= x"C57DFFFC";
end if;
if pc = 53108 then
	inst <= x"8200400C";
end if;
if pc = 53112 then
	inst <= x"07DC0088";
end if;
if pc = 53116 then
	inst <= x"C05C007C";
end if;
if pc = 53120 then
	inst <= x"22640220";
end if;
if pc = 53124 then
	inst <= x"C09C0078";
end if;
if pc = 53128 then
	inst <= x"D4286000";
end if;
if pc = 53132 then
	inst <= x"8200CFC8";
end if;
if pc = 53136 then
	inst <= x"C53C0078";
end if;
if pc = 53140 then
	inst <= x"C4DC007C";
end if;
if pc = 53144 then
	inst <= x"C17DFFFC";
end if;
if pc = 53148 then
	inst <= x"00500000";
end if;
if pc = 53152 then
	inst <= x"00340000";
end if;
if pc = 53156 then
	inst <= x"03DC0088";
end if;
if pc = 53160 then
	inst <= x"037E000C";
end if;
if pc = 53164 then
	inst <= x"C57DFFFC";
end if;
if pc = 53168 then
	inst <= x"82003E98";
end if;
if pc = 53172 then
	inst <= x"07DC0088";
end if;
if pc = 53176 then
	inst <= x"C05C007C";
end if;
if pc = 53180 then
	inst <= x"22640220";
end if;
if pc = 53184 then
	inst <= x"C09C0078";
end if;
if pc = 53188 then
	inst <= x"D4286000";
end if;
if pc = 53192 then
	inst <= x"8200D004";
end if;
if pc = 53196 then
	inst <= x"C53C0078";
end if;
if pc = 53200 then
	inst <= x"C4DC007C";
end if;
if pc = 53204 then
	inst <= x"C17DFFFC";
end if;
if pc = 53208 then
	inst <= x"00500000";
end if;
if pc = 53212 then
	inst <= x"00340000";
end if;
if pc = 53216 then
	inst <= x"03DC0088";
end if;
if pc = 53220 then
	inst <= x"037E000C";
end if;
if pc = 53224 then
	inst <= x"C57DFFFC";
end if;
if pc = 53228 then
	inst <= x"82003CC4";
end if;
if pc = 53232 then
	inst <= x"07DC0088";
end if;
if pc = 53236 then
	inst <= x"C05C007C";
end if;
if pc = 53240 then
	inst <= x"22640220";
end if;
if pc = 53244 then
	inst <= x"C09C0078";
end if;
if pc = 53248 then
	inst <= x"D4286000";
end if;
if pc = 53252 then
	inst <= x"06240001";
end if;
if pc = 53256 then
	inst <= x"8620D100";
end if;
if pc = 53260 then
	inst <= x"22420220";
end if;
if pc = 53264 then
	inst <= x"C07C0074";
end if;
if pc = 53268 then
	inst <= x"D0464000";
end if;
if pc = 53272 then
	inst <= x"C07C0070";
end if;
if pc = 53276 then
	inst <= x"C0860004";
end if;
if pc = 53280 then
	inst <= x"C0A60000";
end if;
if pc = 53284 then
	inst <= x"C0C40004";
end if;
if pc = 53288 then
	inst <= x"02E00001";
end if;
if pc = 53292 then
	inst <= x"82CED0A8";
end if;
if pc = 53296 then
	inst <= x"02E00002";
end if;
if pc = 53300 then
	inst <= x"82CED070";
end if;
if pc = 53304 then
	inst <= x"C49C0080";
end if;
if pc = 53308 then
	inst <= x"C43C0084";
end if;
if pc = 53312 then
	inst <= x"C17DFFFC";
end if;
if pc = 53316 then
	inst <= x"002A0000";
end if;
if pc = 53320 then
	inst <= x"03DC0090";
end if;
if pc = 53324 then
	inst <= x"037E000C";
end if;
if pc = 53328 then
	inst <= x"C57DFFFC";
end if;
if pc = 53332 then
	inst <= x"8200400C";
end if;
if pc = 53336 then
	inst <= x"07DC0090";
end if;
if pc = 53340 then
	inst <= x"C05C0084";
end if;
if pc = 53344 then
	inst <= x"22640220";
end if;
if pc = 53348 then
	inst <= x"C09C0080";
end if;
if pc = 53352 then
	inst <= x"D4286000";
end if;
if pc = 53356 then
	inst <= x"8200D0A4";
end if;
if pc = 53360 then
	inst <= x"C49C0080";
end if;
if pc = 53364 then
	inst <= x"C43C0084";
end if;
if pc = 53368 then
	inst <= x"C17DFFFC";
end if;
if pc = 53372 then
	inst <= x"002A0000";
end if;
if pc = 53376 then
	inst <= x"03DC0090";
end if;
if pc = 53380 then
	inst <= x"037E000C";
end if;
if pc = 53384 then
	inst <= x"C57DFFFC";
end if;
if pc = 53388 then
	inst <= x"82003E98";
end if;
if pc = 53392 then
	inst <= x"07DC0090";
end if;
if pc = 53396 then
	inst <= x"C05C0084";
end if;
if pc = 53400 then
	inst <= x"22640220";
end if;
if pc = 53404 then
	inst <= x"C09C0080";
end if;
if pc = 53408 then
	inst <= x"D4286000";
end if;
if pc = 53412 then
	inst <= x"8200D0DC";
end if;
if pc = 53416 then
	inst <= x"C49C0080";
end if;
if pc = 53420 then
	inst <= x"C43C0084";
end if;
if pc = 53424 then
	inst <= x"C17DFFFC";
end if;
if pc = 53428 then
	inst <= x"002A0000";
end if;
if pc = 53432 then
	inst <= x"03DC0090";
end if;
if pc = 53436 then
	inst <= x"037E000C";
end if;
if pc = 53440 then
	inst <= x"C57DFFFC";
end if;
if pc = 53444 then
	inst <= x"82003CC4";
end if;
if pc = 53448 then
	inst <= x"07DC0090";
end if;
if pc = 53452 then
	inst <= x"C05C0084";
end if;
if pc = 53456 then
	inst <= x"22640220";
end if;
if pc = 53460 then
	inst <= x"C09C0080";
end if;
if pc = 53464 then
	inst <= x"D4286000";
end if;
if pc = 53468 then
	inst <= x"06440001";
end if;
if pc = 53472 then
	inst <= x"C03C0070";
end if;
if pc = 53476 then
	inst <= x"C17DFFFC";
end if;
if pc = 53480 then
	inst <= x"03DC0090";
end if;
if pc = 53484 then
	inst <= x"037E000C";
end if;
if pc = 53488 then
	inst <= x"C57DFFFC";
end if;
if pc = 53492 then
	inst <= x"820042A4";
end if;
if pc = 53496 then
	inst <= x"07DC0090";
end if;
if pc = 53500 then
	inst <= x"8200D100";
end if;
if pc = 53504 then
	inst <= x"8200D104";
end if;
if pc = 53508 then
	inst <= x"C03C006C";
end if;
if pc = 53512 then
	inst <= x"C04201D8";
end if;
if pc = 53516 then
	inst <= x"C07C0008";
end if;
if pc = 53520 then
	inst <= x"C0860000";
end if;
if pc = 53524 then
	inst <= x"06880001";
end if;
if pc = 53528 then
	inst <= x"8680D3D8";
end if;
if pc = 53532 then
	inst <= x"02A000C8";
end if;
if pc = 53536 then
	inst <= x"22C80220";
end if;
if pc = 53540 then
	inst <= x"D0CAC000";
end if;
if pc = 53544 then
	inst <= x"C0E40004";
end if;
if pc = 53548 then
	inst <= x"C1040000";
end if;
if pc = 53552 then
	inst <= x"C12C0004";
end if;
if pc = 53556 then
	inst <= x"03400001";
end if;
if pc = 53560 then
	inst <= x"C45C0088";
end if;
if pc = 53564 then
	inst <= x"C4BC008C";
end if;
if pc = 53568 then
	inst <= x"8334D1C4";
end if;
if pc = 53572 then
	inst <= x"03400002";
end if;
if pc = 53576 then
	inst <= x"8334D188";
end if;
if pc = 53580 then
	inst <= x"C4FC0090";
end if;
if pc = 53584 then
	inst <= x"C49C0094";
end if;
if pc = 53588 then
	inst <= x"C17DFFFC";
end if;
if pc = 53592 then
	inst <= x"004C0000";
end if;
if pc = 53596 then
	inst <= x"00300000";
end if;
if pc = 53600 then
	inst <= x"03DC00A0";
end if;
if pc = 53604 then
	inst <= x"037E000C";
end if;
if pc = 53608 then
	inst <= x"C57DFFFC";
end if;
if pc = 53612 then
	inst <= x"8200400C";
end if;
if pc = 53616 then
	inst <= x"07DC00A0";
end if;
if pc = 53620 then
	inst <= x"C05C0094";
end if;
if pc = 53624 then
	inst <= x"22640220";
end if;
if pc = 53628 then
	inst <= x"C09C0090";
end if;
if pc = 53632 then
	inst <= x"D4286000";
end if;
if pc = 53636 then
	inst <= x"8200D1C0";
end if;
if pc = 53640 then
	inst <= x"C4FC0090";
end if;
if pc = 53644 then
	inst <= x"C49C0094";
end if;
if pc = 53648 then
	inst <= x"C17DFFFC";
end if;
if pc = 53652 then
	inst <= x"004C0000";
end if;
if pc = 53656 then
	inst <= x"00300000";
end if;
if pc = 53660 then
	inst <= x"03DC00A0";
end if;
if pc = 53664 then
	inst <= x"037E000C";
end if;
if pc = 53668 then
	inst <= x"C57DFFFC";
end if;
if pc = 53672 then
	inst <= x"82003E98";
end if;
if pc = 53676 then
	inst <= x"07DC00A0";
end if;
if pc = 53680 then
	inst <= x"C05C0094";
end if;
if pc = 53684 then
	inst <= x"22640220";
end if;
if pc = 53688 then
	inst <= x"C09C0090";
end if;
if pc = 53692 then
	inst <= x"D4286000";
end if;
if pc = 53696 then
	inst <= x"8200D1FC";
end if;
if pc = 53700 then
	inst <= x"C4FC0090";
end if;
if pc = 53704 then
	inst <= x"C49C0094";
end if;
if pc = 53708 then
	inst <= x"C17DFFFC";
end if;
if pc = 53712 then
	inst <= x"004C0000";
end if;
if pc = 53716 then
	inst <= x"00300000";
end if;
if pc = 53720 then
	inst <= x"03DC00A0";
end if;
if pc = 53724 then
	inst <= x"037E000C";
end if;
if pc = 53728 then
	inst <= x"C57DFFFC";
end if;
if pc = 53732 then
	inst <= x"82003CC4";
end if;
if pc = 53736 then
	inst <= x"07DC00A0";
end if;
if pc = 53740 then
	inst <= x"C05C0094";
end if;
if pc = 53744 then
	inst <= x"22640220";
end if;
if pc = 53748 then
	inst <= x"C09C0090";
end if;
if pc = 53752 then
	inst <= x"D4286000";
end if;
if pc = 53756 then
	inst <= x"06240001";
end if;
if pc = 53760 then
	inst <= x"8620D3D4";
end if;
if pc = 53764 then
	inst <= x"22420220";
end if;
if pc = 53768 then
	inst <= x"C07C008C";
end if;
if pc = 53772 then
	inst <= x"D0464000";
end if;
if pc = 53776 then
	inst <= x"C09C0088";
end if;
if pc = 53780 then
	inst <= x"C0A80004";
end if;
if pc = 53784 then
	inst <= x"C0C80000";
end if;
if pc = 53788 then
	inst <= x"C0E40004";
end if;
if pc = 53792 then
	inst <= x"03000001";
end if;
if pc = 53796 then
	inst <= x"82F0D2A0";
end if;
if pc = 53800 then
	inst <= x"03000002";
end if;
if pc = 53804 then
	inst <= x"82F0D268";
end if;
if pc = 53808 then
	inst <= x"C4BC0098";
end if;
if pc = 53812 then
	inst <= x"C43C009C";
end if;
if pc = 53816 then
	inst <= x"C17DFFFC";
end if;
if pc = 53820 then
	inst <= x"002C0000";
end if;
if pc = 53824 then
	inst <= x"03DC00A8";
end if;
if pc = 53828 then
	inst <= x"037E000C";
end if;
if pc = 53832 then
	inst <= x"C57DFFFC";
end if;
if pc = 53836 then
	inst <= x"8200400C";
end if;
if pc = 53840 then
	inst <= x"07DC00A8";
end if;
if pc = 53844 then
	inst <= x"C05C009C";
end if;
if pc = 53848 then
	inst <= x"22640220";
end if;
if pc = 53852 then
	inst <= x"C09C0098";
end if;
if pc = 53856 then
	inst <= x"D4286000";
end if;
if pc = 53860 then
	inst <= x"8200D29C";
end if;
if pc = 53864 then
	inst <= x"C4BC0098";
end if;
if pc = 53868 then
	inst <= x"C43C009C";
end if;
if pc = 53872 then
	inst <= x"C17DFFFC";
end if;
if pc = 53876 then
	inst <= x"002C0000";
end if;
if pc = 53880 then
	inst <= x"03DC00A8";
end if;
if pc = 53884 then
	inst <= x"037E000C";
end if;
if pc = 53888 then
	inst <= x"C57DFFFC";
end if;
if pc = 53892 then
	inst <= x"82003E98";
end if;
if pc = 53896 then
	inst <= x"07DC00A8";
end if;
if pc = 53900 then
	inst <= x"C05C009C";
end if;
if pc = 53904 then
	inst <= x"22640220";
end if;
if pc = 53908 then
	inst <= x"C09C0098";
end if;
if pc = 53912 then
	inst <= x"D4286000";
end if;
if pc = 53916 then
	inst <= x"8200D2D4";
end if;
if pc = 53920 then
	inst <= x"C4BC0098";
end if;
if pc = 53924 then
	inst <= x"C43C009C";
end if;
if pc = 53928 then
	inst <= x"C17DFFFC";
end if;
if pc = 53932 then
	inst <= x"002C0000";
end if;
if pc = 53936 then
	inst <= x"03DC00A8";
end if;
if pc = 53940 then
	inst <= x"037E000C";
end if;
if pc = 53944 then
	inst <= x"C57DFFFC";
end if;
if pc = 53948 then
	inst <= x"82003CC4";
end if;
if pc = 53952 then
	inst <= x"07DC00A8";
end if;
if pc = 53956 then
	inst <= x"C05C009C";
end if;
if pc = 53960 then
	inst <= x"22640220";
end if;
if pc = 53964 then
	inst <= x"C09C0098";
end if;
if pc = 53968 then
	inst <= x"D4286000";
end if;
if pc = 53972 then
	inst <= x"06240001";
end if;
if pc = 53976 then
	inst <= x"8620D3D0";
end if;
if pc = 53980 then
	inst <= x"22420220";
end if;
if pc = 53984 then
	inst <= x"C07C008C";
end if;
if pc = 53988 then
	inst <= x"D0464000";
end if;
if pc = 53992 then
	inst <= x"C07C0088";
end if;
if pc = 53996 then
	inst <= x"C0860004";
end if;
if pc = 54000 then
	inst <= x"C0A60000";
end if;
if pc = 54004 then
	inst <= x"C0C40004";
end if;
if pc = 54008 then
	inst <= x"02E00001";
end if;
if pc = 54012 then
	inst <= x"82CED378";
end if;
if pc = 54016 then
	inst <= x"02E00002";
end if;
if pc = 54020 then
	inst <= x"82CED340";
end if;
if pc = 54024 then
	inst <= x"C49C00A0";
end if;
if pc = 54028 then
	inst <= x"C43C00A4";
end if;
if pc = 54032 then
	inst <= x"C17DFFFC";
end if;
if pc = 54036 then
	inst <= x"002A0000";
end if;
if pc = 54040 then
	inst <= x"03DC00B0";
end if;
if pc = 54044 then
	inst <= x"037E000C";
end if;
if pc = 54048 then
	inst <= x"C57DFFFC";
end if;
if pc = 54052 then
	inst <= x"8200400C";
end if;
if pc = 54056 then
	inst <= x"07DC00B0";
end if;
if pc = 54060 then
	inst <= x"C05C00A4";
end if;
if pc = 54064 then
	inst <= x"22640220";
end if;
if pc = 54068 then
	inst <= x"C09C00A0";
end if;
if pc = 54072 then
	inst <= x"D4286000";
end if;
if pc = 54076 then
	inst <= x"8200D374";
end if;
if pc = 54080 then
	inst <= x"C49C00A0";
end if;
if pc = 54084 then
	inst <= x"C43C00A4";
end if;
if pc = 54088 then
	inst <= x"C17DFFFC";
end if;
if pc = 54092 then
	inst <= x"002A0000";
end if;
if pc = 54096 then
	inst <= x"03DC00B0";
end if;
if pc = 54100 then
	inst <= x"037E000C";
end if;
if pc = 54104 then
	inst <= x"C57DFFFC";
end if;
if pc = 54108 then
	inst <= x"82003E98";
end if;
if pc = 54112 then
	inst <= x"07DC00B0";
end if;
if pc = 54116 then
	inst <= x"C05C00A4";
end if;
if pc = 54120 then
	inst <= x"22640220";
end if;
if pc = 54124 then
	inst <= x"C09C00A0";
end if;
if pc = 54128 then
	inst <= x"D4286000";
end if;
if pc = 54132 then
	inst <= x"8200D3AC";
end if;
if pc = 54136 then
	inst <= x"C49C00A0";
end if;
if pc = 54140 then
	inst <= x"C43C00A4";
end if;
if pc = 54144 then
	inst <= x"C17DFFFC";
end if;
if pc = 54148 then
	inst <= x"002A0000";
end if;
if pc = 54152 then
	inst <= x"03DC00B0";
end if;
if pc = 54156 then
	inst <= x"037E000C";
end if;
if pc = 54160 then
	inst <= x"C57DFFFC";
end if;
if pc = 54164 then
	inst <= x"82003CC4";
end if;
if pc = 54168 then
	inst <= x"07DC00B0";
end if;
if pc = 54172 then
	inst <= x"C05C00A4";
end if;
if pc = 54176 then
	inst <= x"22640220";
end if;
if pc = 54180 then
	inst <= x"C09C00A0";
end if;
if pc = 54184 then
	inst <= x"D4286000";
end if;
if pc = 54188 then
	inst <= x"06440001";
end if;
if pc = 54192 then
	inst <= x"C03C0088";
end if;
if pc = 54196 then
	inst <= x"C17DFFFC";
end if;
if pc = 54200 then
	inst <= x"03DC00B0";
end if;
if pc = 54204 then
	inst <= x"037E000C";
end if;
if pc = 54208 then
	inst <= x"C57DFFFC";
end if;
if pc = 54212 then
	inst <= x"820042A4";
end if;
if pc = 54216 then
	inst <= x"07DC00B0";
end if;
if pc = 54220 then
	inst <= x"8200D3D0";
end if;
if pc = 54224 then
	inst <= x"8200D3D4";
end if;
if pc = 54228 then
	inst <= x"8200D3D8";
end if;
if pc = 54232 then
	inst <= x"02400075";
end if;
if pc = 54236 then
	inst <= x"C03C006C";
end if;
if pc = 54240 then
	inst <= x"C17DFFFC";
end if;
if pc = 54244 then
	inst <= x"03DC00B0";
end if;
if pc = 54248 then
	inst <= x"037E000C";
end if;
if pc = 54252 then
	inst <= x"C57DFFFC";
end if;
if pc = 54256 then
	inst <= x"8200BD10";
end if;
if pc = 54260 then
	inst <= x"07DC00B0";
end if;
if pc = 54264 then
	inst <= x"C03C0068";
end if;
if pc = 54268 then
	inst <= x"06220001";
end if;
if pc = 54272 then
	inst <= x"8620D758";
end if;
if pc = 54276 then
	inst <= x"22420220";
end if;
if pc = 54280 then
	inst <= x"C07C0000";
end if;
if pc = 54284 then
	inst <= x"D0464000";
end if;
if pc = 54288 then
	inst <= x"C08401DC";
end if;
if pc = 54292 then
	inst <= x"C0BC0008";
end if;
if pc = 54296 then
	inst <= x"C0AA0000";
end if;
if pc = 54300 then
	inst <= x"06AA0001";
end if;
if pc = 54304 then
	inst <= x"C43C00A8";
end if;
if pc = 54308 then
	inst <= x"C45C00AC";
end if;
if pc = 54312 then
	inst <= x"86A0D6E8";
end if;
if pc = 54316 then
	inst <= x"02C000C8";
end if;
if pc = 54320 then
	inst <= x"22EA0220";
end if;
if pc = 54324 then
	inst <= x"D0ECE000";
end if;
if pc = 54328 then
	inst <= x"C1080004";
end if;
if pc = 54332 then
	inst <= x"C1280000";
end if;
if pc = 54336 then
	inst <= x"C14E0004";
end if;
if pc = 54340 then
	inst <= x"02600001";
end if;
if pc = 54344 then
	inst <= x"C49C00B0";
end if;
if pc = 54348 then
	inst <= x"C4DC00B4";
end if;
if pc = 54352 then
	inst <= x"8346D4D4";
end if;
if pc = 54356 then
	inst <= x"02600002";
end if;
if pc = 54360 then
	inst <= x"8346D498";
end if;
if pc = 54364 then
	inst <= x"C51C00B8";
end if;
if pc = 54368 then
	inst <= x"C4BC00BC";
end if;
if pc = 54372 then
	inst <= x"C17DFFFC";
end if;
if pc = 54376 then
	inst <= x"004E0000";
end if;
if pc = 54380 then
	inst <= x"00320000";
end if;
if pc = 54384 then
	inst <= x"03DC00C8";
end if;
if pc = 54388 then
	inst <= x"037E000C";
end if;
if pc = 54392 then
	inst <= x"C57DFFFC";
end if;
if pc = 54396 then
	inst <= x"8200400C";
end if;
if pc = 54400 then
	inst <= x"07DC00C8";
end if;
if pc = 54404 then
	inst <= x"C05C00BC";
end if;
if pc = 54408 then
	inst <= x"22640220";
end if;
if pc = 54412 then
	inst <= x"C09C00B8";
end if;
if pc = 54416 then
	inst <= x"D4286000";
end if;
if pc = 54420 then
	inst <= x"8200D4D0";
end if;
if pc = 54424 then
	inst <= x"C51C00B8";
end if;
if pc = 54428 then
	inst <= x"C4BC00BC";
end if;
if pc = 54432 then
	inst <= x"C17DFFFC";
end if;
if pc = 54436 then
	inst <= x"004E0000";
end if;
if pc = 54440 then
	inst <= x"00320000";
end if;
if pc = 54444 then
	inst <= x"03DC00C8";
end if;
if pc = 54448 then
	inst <= x"037E000C";
end if;
if pc = 54452 then
	inst <= x"C57DFFFC";
end if;
if pc = 54456 then
	inst <= x"82003E98";
end if;
if pc = 54460 then
	inst <= x"07DC00C8";
end if;
if pc = 54464 then
	inst <= x"C05C00BC";
end if;
if pc = 54468 then
	inst <= x"22640220";
end if;
if pc = 54472 then
	inst <= x"C09C00B8";
end if;
if pc = 54476 then
	inst <= x"D4286000";
end if;
if pc = 54480 then
	inst <= x"8200D50C";
end if;
if pc = 54484 then
	inst <= x"C51C00B8";
end if;
if pc = 54488 then
	inst <= x"C4BC00BC";
end if;
if pc = 54492 then
	inst <= x"C17DFFFC";
end if;
if pc = 54496 then
	inst <= x"004E0000";
end if;
if pc = 54500 then
	inst <= x"00320000";
end if;
if pc = 54504 then
	inst <= x"03DC00C8";
end if;
if pc = 54508 then
	inst <= x"037E000C";
end if;
if pc = 54512 then
	inst <= x"C57DFFFC";
end if;
if pc = 54516 then
	inst <= x"82003CC4";
end if;
if pc = 54520 then
	inst <= x"07DC00C8";
end if;
if pc = 54524 then
	inst <= x"C05C00BC";
end if;
if pc = 54528 then
	inst <= x"22640220";
end if;
if pc = 54532 then
	inst <= x"C09C00B8";
end if;
if pc = 54536 then
	inst <= x"D4286000";
end if;
if pc = 54540 then
	inst <= x"06240001";
end if;
if pc = 54544 then
	inst <= x"8620D6E4";
end if;
if pc = 54548 then
	inst <= x"22420220";
end if;
if pc = 54552 then
	inst <= x"C07C00B4";
end if;
if pc = 54556 then
	inst <= x"D0464000";
end if;
if pc = 54560 then
	inst <= x"C09C00B0";
end if;
if pc = 54564 then
	inst <= x"C0A80004";
end if;
if pc = 54568 then
	inst <= x"C0C80000";
end if;
if pc = 54572 then
	inst <= x"C0E40004";
end if;
if pc = 54576 then
	inst <= x"03000001";
end if;
if pc = 54580 then
	inst <= x"82F0D5B0";
end if;
if pc = 54584 then
	inst <= x"03000002";
end if;
if pc = 54588 then
	inst <= x"82F0D578";
end if;
if pc = 54592 then
	inst <= x"C4BC00C0";
end if;
if pc = 54596 then
	inst <= x"C43C00C4";
end if;
if pc = 54600 then
	inst <= x"C17DFFFC";
end if;
if pc = 54604 then
	inst <= x"002C0000";
end if;
if pc = 54608 then
	inst <= x"03DC00D0";
end if;
if pc = 54612 then
	inst <= x"037E000C";
end if;
if pc = 54616 then
	inst <= x"C57DFFFC";
end if;
if pc = 54620 then
	inst <= x"8200400C";
end if;
if pc = 54624 then
	inst <= x"07DC00D0";
end if;
if pc = 54628 then
	inst <= x"C05C00C4";
end if;
if pc = 54632 then
	inst <= x"22640220";
end if;
if pc = 54636 then
	inst <= x"C09C00C0";
end if;
if pc = 54640 then
	inst <= x"D4286000";
end if;
if pc = 54644 then
	inst <= x"8200D5AC";
end if;
if pc = 54648 then
	inst <= x"C4BC00C0";
end if;
if pc = 54652 then
	inst <= x"C43C00C4";
end if;
if pc = 54656 then
	inst <= x"C17DFFFC";
end if;
if pc = 54660 then
	inst <= x"002C0000";
end if;
if pc = 54664 then
	inst <= x"03DC00D0";
end if;
if pc = 54668 then
	inst <= x"037E000C";
end if;
if pc = 54672 then
	inst <= x"C57DFFFC";
end if;
if pc = 54676 then
	inst <= x"82003E98";
end if;
if pc = 54680 then
	inst <= x"07DC00D0";
end if;
if pc = 54684 then
	inst <= x"C05C00C4";
end if;
if pc = 54688 then
	inst <= x"22640220";
end if;
if pc = 54692 then
	inst <= x"C09C00C0";
end if;
if pc = 54696 then
	inst <= x"D4286000";
end if;
if pc = 54700 then
	inst <= x"8200D5E4";
end if;
if pc = 54704 then
	inst <= x"C4BC00C0";
end if;
if pc = 54708 then
	inst <= x"C43C00C4";
end if;
if pc = 54712 then
	inst <= x"C17DFFFC";
end if;
if pc = 54716 then
	inst <= x"002C0000";
end if;
if pc = 54720 then
	inst <= x"03DC00D0";
end if;
if pc = 54724 then
	inst <= x"037E000C";
end if;
if pc = 54728 then
	inst <= x"C57DFFFC";
end if;
if pc = 54732 then
	inst <= x"82003CC4";
end if;
if pc = 54736 then
	inst <= x"07DC00D0";
end if;
if pc = 54740 then
	inst <= x"C05C00C4";
end if;
if pc = 54744 then
	inst <= x"22640220";
end if;
if pc = 54748 then
	inst <= x"C09C00C0";
end if;
if pc = 54752 then
	inst <= x"D4286000";
end if;
if pc = 54756 then
	inst <= x"06240001";
end if;
if pc = 54760 then
	inst <= x"8620D6E0";
end if;
if pc = 54764 then
	inst <= x"22420220";
end if;
if pc = 54768 then
	inst <= x"C07C00B4";
end if;
if pc = 54772 then
	inst <= x"D0464000";
end if;
if pc = 54776 then
	inst <= x"C07C00B0";
end if;
if pc = 54780 then
	inst <= x"C0860004";
end if;
if pc = 54784 then
	inst <= x"C0A60000";
end if;
if pc = 54788 then
	inst <= x"C0C40004";
end if;
if pc = 54792 then
	inst <= x"02E00001";
end if;
if pc = 54796 then
	inst <= x"82CED688";
end if;
if pc = 54800 then
	inst <= x"02E00002";
end if;
if pc = 54804 then
	inst <= x"82CED650";
end if;
if pc = 54808 then
	inst <= x"C49C00C8";
end if;
if pc = 54812 then
	inst <= x"C43C00CC";
end if;
if pc = 54816 then
	inst <= x"C17DFFFC";
end if;
if pc = 54820 then
	inst <= x"002A0000";
end if;
if pc = 54824 then
	inst <= x"03DC00D8";
end if;
if pc = 54828 then
	inst <= x"037E000C";
end if;
if pc = 54832 then
	inst <= x"C57DFFFC";
end if;
if pc = 54836 then
	inst <= x"8200400C";
end if;
if pc = 54840 then
	inst <= x"07DC00D8";
end if;
if pc = 54844 then
	inst <= x"C05C00CC";
end if;
if pc = 54848 then
	inst <= x"22640220";
end if;
if pc = 54852 then
	inst <= x"C09C00C8";
end if;
if pc = 54856 then
	inst <= x"D4286000";
end if;
if pc = 54860 then
	inst <= x"8200D684";
end if;
if pc = 54864 then
	inst <= x"C49C00C8";
end if;
if pc = 54868 then
	inst <= x"C43C00CC";
end if;
if pc = 54872 then
	inst <= x"C17DFFFC";
end if;
if pc = 54876 then
	inst <= x"002A0000";
end if;
if pc = 54880 then
	inst <= x"03DC00D8";
end if;
if pc = 54884 then
	inst <= x"037E000C";
end if;
if pc = 54888 then
	inst <= x"C57DFFFC";
end if;
if pc = 54892 then
	inst <= x"82003E98";
end if;
if pc = 54896 then
	inst <= x"07DC00D8";
end if;
if pc = 54900 then
	inst <= x"C05C00CC";
end if;
if pc = 54904 then
	inst <= x"22640220";
end if;
if pc = 54908 then
	inst <= x"C09C00C8";
end if;
if pc = 54912 then
	inst <= x"D4286000";
end if;
if pc = 54916 then
	inst <= x"8200D6BC";
end if;
if pc = 54920 then
	inst <= x"C49C00C8";
end if;
if pc = 54924 then
	inst <= x"C43C00CC";
end if;
if pc = 54928 then
	inst <= x"C17DFFFC";
end if;
if pc = 54932 then
	inst <= x"002A0000";
end if;
if pc = 54936 then
	inst <= x"03DC00D8";
end if;
if pc = 54940 then
	inst <= x"037E000C";
end if;
if pc = 54944 then
	inst <= x"C57DFFFC";
end if;
if pc = 54948 then
	inst <= x"82003CC4";
end if;
if pc = 54952 then
	inst <= x"07DC00D8";
end if;
if pc = 54956 then
	inst <= x"C05C00CC";
end if;
if pc = 54960 then
	inst <= x"22640220";
end if;
if pc = 54964 then
	inst <= x"C09C00C8";
end if;
if pc = 54968 then
	inst <= x"D4286000";
end if;
if pc = 54972 then
	inst <= x"06440001";
end if;
if pc = 54976 then
	inst <= x"C03C00B0";
end if;
if pc = 54980 then
	inst <= x"C17DFFFC";
end if;
if pc = 54984 then
	inst <= x"03DC00D8";
end if;
if pc = 54988 then
	inst <= x"037E000C";
end if;
if pc = 54992 then
	inst <= x"C57DFFFC";
end if;
if pc = 54996 then
	inst <= x"820042A4";
end if;
if pc = 55000 then
	inst <= x"07DC00D8";
end if;
if pc = 55004 then
	inst <= x"8200D6E0";
end if;
if pc = 55008 then
	inst <= x"8200D6E4";
end if;
if pc = 55012 then
	inst <= x"8200D6E8";
end if;
if pc = 55016 then
	inst <= x"02400076";
end if;
if pc = 55020 then
	inst <= x"C03C00AC";
end if;
if pc = 55024 then
	inst <= x"C17DFFFC";
end if;
if pc = 55028 then
	inst <= x"03DC00D8";
end if;
if pc = 55032 then
	inst <= x"037E000C";
end if;
if pc = 55036 then
	inst <= x"C57DFFFC";
end if;
if pc = 55040 then
	inst <= x"8200BD10";
end if;
if pc = 55044 then
	inst <= x"07DC00D8";
end if;
if pc = 55048 then
	inst <= x"C03C00A8";
end if;
if pc = 55052 then
	inst <= x"06220001";
end if;
if pc = 55056 then
	inst <= x"8620D754";
end if;
if pc = 55060 then
	inst <= x"22420220";
end if;
if pc = 55064 then
	inst <= x"C07C0000";
end if;
if pc = 55068 then
	inst <= x"D0464000";
end if;
if pc = 55072 then
	inst <= x"02600077";
end if;
if pc = 55076 then
	inst <= x"C43C00D0";
end if;
if pc = 55080 then
	inst <= x"C17DFFFC";
end if;
if pc = 55084 then
	inst <= x"00240000";
end if;
if pc = 55088 then
	inst <= x"00460000";
end if;
if pc = 55092 then
	inst <= x"03DC00DC";
end if;
if pc = 55096 then
	inst <= x"037E000C";
end if;
if pc = 55100 then
	inst <= x"C57DFFFC";
end if;
if pc = 55104 then
	inst <= x"8200BD10";
end if;
if pc = 55108 then
	inst <= x"07DC00DC";
end if;
if pc = 55112 then
	inst <= x"C03C00D0";
end if;
if pc = 55116 then
	inst <= x"06220001";
end if;
if pc = 55120 then
	inst <= x"8200C714";
end if;
if pc = 55124 then
	inst <= x"C1FDFFFC";
end if;
if pc = 55128 then
	inst <= x"C1FDFFFC";
end if;
if pc = 55132 then
	inst <= x"C1FDFFFC";
end if;
if pc = 55136 then
	inst <= x"C1FDFFFC";
end if;
if pc = 55140 then
	inst <= x"22220220";
end if;
if pc = 55144 then
	inst <= x"02600640";
end if;
if pc = 55148 then
	inst <= x"C0860000";
end if;
if pc = 55152 then
	inst <= x"C82000A8";
end if;
if pc = 55156 then
	inst <= x"C044001C";
end if;
if pc = 55160 then
	inst <= x"C8440000";
end if;
if pc = 55164 then
	inst <= x"44224000";
end if;
if pc = 55168 then
	inst <= x"024001D0";
end if;
if pc = 55172 then
	inst <= x"C8440000";
end if;
if pc = 55176 then
	inst <= x"44404000";
end if;
if pc = 55180 then
	inst <= x"C8640004";
end if;
if pc = 55184 then
	inst <= x"44606000";
end if;
if pc = 55188 then
	inst <= x"C8840008";
end if;
if pc = 55192 then
	inst <= x"44808000";
end if;
if pc = 55196 then
	inst <= x"02A20001";
end if;
if pc = 55200 then
	inst <= x"C8A40000";
end if;
if pc = 55204 then
	inst <= x"02C00003";
end if;
if pc = 55208 then
	inst <= x"40C00000";
end if;
if pc = 55212 then
	inst <= x"C47C0000";
end if;
if pc = 55216 then
	inst <= x"CC5C0008";
end if;
if pc = 55220 then
	inst <= x"CCDC0010";
end if;
if pc = 55224 then
	inst <= x"C45C0018";
end if;
if pc = 55228 then
	inst <= x"C43C001C";
end if;
if pc = 55232 then
	inst <= x"C49C0020";
end if;
if pc = 55236 then
	inst <= x"C4BC0024";
end if;
if pc = 55240 then
	inst <= x"CC3C0028";
end if;
if pc = 55244 then
	inst <= x"CC9C0030";
end if;
if pc = 55248 then
	inst <= x"CC7C0038";
end if;
if pc = 55252 then
	inst <= x"CCBC0040";
end if;
if pc = 55256 then
	inst <= x"C17DFFFC";
end if;
if pc = 55260 then
	inst <= x"002C0000";
end if;
if pc = 55264 then
	inst <= x"4020C000";
end if;
if pc = 55268 then
	inst <= x"03DC0050";
end if;
if pc = 55272 then
	inst <= x"037E000C";
end if;
if pc = 55276 then
	inst <= x"C57DFFFC";
end if;
if pc = 55280 then
	inst <= x"8200081C";
end if;
if pc = 55284 then
	inst <= x"07DC0050";
end if;
if pc = 55288 then
	inst <= x"00420000";
end if;
if pc = 55292 then
	inst <= x"022000C4";
end if;
if pc = 55296 then
	inst <= x"C0620000";
end if;
if pc = 55300 then
	inst <= x"C43C0048";
end if;
if pc = 55304 then
	inst <= x"C45C004C";
end if;
if pc = 55308 then
	inst <= x"C17DFFFC";
end if;
if pc = 55312 then
	inst <= x"00260000";
end if;
if pc = 55316 then
	inst <= x"03DC0058";
end if;
if pc = 55320 then
	inst <= x"037E000C";
end if;
if pc = 55324 then
	inst <= x"C57DFFFC";
end if;
if pc = 55328 then
	inst <= x"8200081C";
end if;
if pc = 55332 then
	inst <= x"07DC0058";
end if;
if pc = 55336 then
	inst <= x"005A0000";
end if;
if pc = 55340 then
	inst <= x"03BA0008";
end if;
if pc = 55344 then
	inst <= x"C4240004";
end if;
if pc = 55348 then
	inst <= x"C07C004C";
end if;
if pc = 55352 then
	inst <= x"C4640000";
end if;
if pc = 55356 then
	inst <= x"C83C0040";
end if;
if pc = 55360 then
	inst <= x"CC260000";
end if;
if pc = 55364 then
	inst <= x"C83C0038";
end if;
if pc = 55368 then
	inst <= x"CC260004";
end if;
if pc = 55372 then
	inst <= x"C85C0030";
end if;
if pc = 55376 then
	inst <= x"CC460008";
end if;
if pc = 55380 then
	inst <= x"C09C0048";
end if;
if pc = 55384 then
	inst <= x"C0A80000";
end if;
if pc = 55388 then
	inst <= x"06AA0001";
end if;
if pc = 55392 then
	inst <= x"C45C0050";
end if;
if pc = 55396 then
	inst <= x"86A0DB00";
end if;
if pc = 55400 then
	inst <= x"02C000C8";
end if;
if pc = 55404 then
	inst <= x"22EA0220";
end if;
if pc = 55408 then
	inst <= x"D0ECE000";
end if;
if pc = 55412 then
	inst <= x"C10E0004";
end if;
if pc = 55416 then
	inst <= x"03200001";
end if;
if pc = 55420 then
	inst <= x"C4DC0054";
end if;
if pc = 55424 then
	inst <= x"8312D904";
end if;
if pc = 55428 then
	inst <= x"03200002";
end if;
if pc = 55432 then
	inst <= x"8312D8C8";
end if;
if pc = 55436 then
	inst <= x"C43C0058";
end if;
if pc = 55440 then
	inst <= x"C4BC005C";
end if;
if pc = 55444 then
	inst <= x"C17DFFFC";
end if;
if pc = 55448 then
	inst <= x"004E0000";
end if;
if pc = 55452 then
	inst <= x"00260000";
end if;
if pc = 55456 then
	inst <= x"03DC0068";
end if;
if pc = 55460 then
	inst <= x"037E000C";
end if;
if pc = 55464 then
	inst <= x"C57DFFFC";
end if;
if pc = 55468 then
	inst <= x"8200400C";
end if;
if pc = 55472 then
	inst <= x"07DC0068";
end if;
if pc = 55476 then
	inst <= x"C05C005C";
end if;
if pc = 55480 then
	inst <= x"22640220";
end if;
if pc = 55484 then
	inst <= x"C09C0058";
end if;
if pc = 55488 then
	inst <= x"D4286000";
end if;
if pc = 55492 then
	inst <= x"8200D900";
end if;
if pc = 55496 then
	inst <= x"C43C0058";
end if;
if pc = 55500 then
	inst <= x"C4BC005C";
end if;
if pc = 55504 then
	inst <= x"C17DFFFC";
end if;
if pc = 55508 then
	inst <= x"004E0000";
end if;
if pc = 55512 then
	inst <= x"00260000";
end if;
if pc = 55516 then
	inst <= x"03DC0068";
end if;
if pc = 55520 then
	inst <= x"037E000C";
end if;
if pc = 55524 then
	inst <= x"C57DFFFC";
end if;
if pc = 55528 then
	inst <= x"82003E98";
end if;
if pc = 55532 then
	inst <= x"07DC0068";
end if;
if pc = 55536 then
	inst <= x"C05C005C";
end if;
if pc = 55540 then
	inst <= x"22640220";
end if;
if pc = 55544 then
	inst <= x"C09C0058";
end if;
if pc = 55548 then
	inst <= x"D4286000";
end if;
if pc = 55552 then
	inst <= x"8200D93C";
end if;
if pc = 55556 then
	inst <= x"C43C0058";
end if;
if pc = 55560 then
	inst <= x"C4BC005C";
end if;
if pc = 55564 then
	inst <= x"C17DFFFC";
end if;
if pc = 55568 then
	inst <= x"004E0000";
end if;
if pc = 55572 then
	inst <= x"00260000";
end if;
if pc = 55576 then
	inst <= x"03DC0068";
end if;
if pc = 55580 then
	inst <= x"037E000C";
end if;
if pc = 55584 then
	inst <= x"C57DFFFC";
end if;
if pc = 55588 then
	inst <= x"82003CC4";
end if;
if pc = 55592 then
	inst <= x"07DC0068";
end if;
if pc = 55596 then
	inst <= x"C05C005C";
end if;
if pc = 55600 then
	inst <= x"22640220";
end if;
if pc = 55604 then
	inst <= x"C09C0058";
end if;
if pc = 55608 then
	inst <= x"D4286000";
end if;
if pc = 55612 then
	inst <= x"06240001";
end if;
if pc = 55616 then
	inst <= x"8620DAFC";
end if;
if pc = 55620 then
	inst <= x"22420220";
end if;
if pc = 55624 then
	inst <= x"C07C0054";
end if;
if pc = 55628 then
	inst <= x"D0464000";
end if;
if pc = 55632 then
	inst <= x"C0A40004";
end if;
if pc = 55636 then
	inst <= x"02C00001";
end if;
if pc = 55640 then
	inst <= x"82ACD9D4";
end if;
if pc = 55644 then
	inst <= x"02C00002";
end if;
if pc = 55648 then
	inst <= x"82ACD99C";
end if;
if pc = 55652 then
	inst <= x"C0BC004C";
end if;
if pc = 55656 then
	inst <= x"C43C0060";
end if;
if pc = 55660 then
	inst <= x"C17DFFFC";
end if;
if pc = 55664 then
	inst <= x"002A0000";
end if;
if pc = 55668 then
	inst <= x"03DC006C";
end if;
if pc = 55672 then
	inst <= x"037E000C";
end if;
if pc = 55676 then
	inst <= x"C57DFFFC";
end if;
if pc = 55680 then
	inst <= x"8200400C";
end if;
if pc = 55684 then
	inst <= x"07DC006C";
end if;
if pc = 55688 then
	inst <= x"C05C0060";
end if;
if pc = 55692 then
	inst <= x"22640220";
end if;
if pc = 55696 then
	inst <= x"C09C0058";
end if;
if pc = 55700 then
	inst <= x"D4286000";
end if;
if pc = 55704 then
	inst <= x"8200D9D0";
end if;
if pc = 55708 then
	inst <= x"C0BC004C";
end if;
if pc = 55712 then
	inst <= x"C43C0060";
end if;
if pc = 55716 then
	inst <= x"C17DFFFC";
end if;
if pc = 55720 then
	inst <= x"002A0000";
end if;
if pc = 55724 then
	inst <= x"03DC006C";
end if;
if pc = 55728 then
	inst <= x"037E000C";
end if;
if pc = 55732 then
	inst <= x"C57DFFFC";
end if;
if pc = 55736 then
	inst <= x"82003E98";
end if;
if pc = 55740 then
	inst <= x"07DC006C";
end if;
if pc = 55744 then
	inst <= x"C05C0060";
end if;
if pc = 55748 then
	inst <= x"22640220";
end if;
if pc = 55752 then
	inst <= x"C09C0058";
end if;
if pc = 55756 then
	inst <= x"D4286000";
end if;
if pc = 55760 then
	inst <= x"8200DA08";
end if;
if pc = 55764 then
	inst <= x"C0BC004C";
end if;
if pc = 55768 then
	inst <= x"C43C0060";
end if;
if pc = 55772 then
	inst <= x"C17DFFFC";
end if;
if pc = 55776 then
	inst <= x"002A0000";
end if;
if pc = 55780 then
	inst <= x"03DC006C";
end if;
if pc = 55784 then
	inst <= x"037E000C";
end if;
if pc = 55788 then
	inst <= x"C57DFFFC";
end if;
if pc = 55792 then
	inst <= x"82003CC4";
end if;
if pc = 55796 then
	inst <= x"07DC006C";
end if;
if pc = 55800 then
	inst <= x"C05C0060";
end if;
if pc = 55804 then
	inst <= x"22640220";
end if;
if pc = 55808 then
	inst <= x"C09C0058";
end if;
if pc = 55812 then
	inst <= x"D4286000";
end if;
if pc = 55816 then
	inst <= x"06240001";
end if;
if pc = 55820 then
	inst <= x"8620DAF8";
end if;
if pc = 55824 then
	inst <= x"22420220";
end if;
if pc = 55828 then
	inst <= x"C07C0054";
end if;
if pc = 55832 then
	inst <= x"D0464000";
end if;
if pc = 55836 then
	inst <= x"C0640004";
end if;
if pc = 55840 then
	inst <= x"02A00001";
end if;
if pc = 55844 then
	inst <= x"826ADAA0";
end if;
if pc = 55848 then
	inst <= x"02A00002";
end if;
if pc = 55852 then
	inst <= x"826ADA68";
end if;
if pc = 55856 then
	inst <= x"C07C004C";
end if;
if pc = 55860 then
	inst <= x"C43C0064";
end if;
if pc = 55864 then
	inst <= x"C17DFFFC";
end if;
if pc = 55868 then
	inst <= x"00260000";
end if;
if pc = 55872 then
	inst <= x"03DC0070";
end if;
if pc = 55876 then
	inst <= x"037E000C";
end if;
if pc = 55880 then
	inst <= x"C57DFFFC";
end if;
if pc = 55884 then
	inst <= x"8200400C";
end if;
if pc = 55888 then
	inst <= x"07DC0070";
end if;
if pc = 55892 then
	inst <= x"C05C0064";
end if;
if pc = 55896 then
	inst <= x"22640220";
end if;
if pc = 55900 then
	inst <= x"C09C0058";
end if;
if pc = 55904 then
	inst <= x"D4286000";
end if;
if pc = 55908 then
	inst <= x"8200DA9C";
end if;
if pc = 55912 then
	inst <= x"C07C004C";
end if;
if pc = 55916 then
	inst <= x"C43C0064";
end if;
if pc = 55920 then
	inst <= x"C17DFFFC";
end if;
if pc = 55924 then
	inst <= x"00260000";
end if;
if pc = 55928 then
	inst <= x"03DC0070";
end if;
if pc = 55932 then
	inst <= x"037E000C";
end if;
if pc = 55936 then
	inst <= x"C57DFFFC";
end if;
if pc = 55940 then
	inst <= x"82003E98";
end if;
if pc = 55944 then
	inst <= x"07DC0070";
end if;
if pc = 55948 then
	inst <= x"C05C0064";
end if;
if pc = 55952 then
	inst <= x"22640220";
end if;
if pc = 55956 then
	inst <= x"C09C0058";
end if;
if pc = 55960 then
	inst <= x"D4286000";
end if;
if pc = 55964 then
	inst <= x"8200DAD4";
end if;
if pc = 55968 then
	inst <= x"C07C004C";
end if;
if pc = 55972 then
	inst <= x"C43C0064";
end if;
if pc = 55976 then
	inst <= x"C17DFFFC";
end if;
if pc = 55980 then
	inst <= x"00260000";
end if;
if pc = 55984 then
	inst <= x"03DC0070";
end if;
if pc = 55988 then
	inst <= x"037E000C";
end if;
if pc = 55992 then
	inst <= x"C57DFFFC";
end if;
if pc = 55996 then
	inst <= x"82003CC4";
end if;
if pc = 56000 then
	inst <= x"07DC0070";
end if;
if pc = 56004 then
	inst <= x"C05C0064";
end if;
if pc = 56008 then
	inst <= x"22640220";
end if;
if pc = 56012 then
	inst <= x"C09C0058";
end if;
if pc = 56016 then
	inst <= x"D4286000";
end if;
if pc = 56020 then
	inst <= x"06440001";
end if;
if pc = 56024 then
	inst <= x"C03C0050";
end if;
if pc = 56028 then
	inst <= x"C17DFFFC";
end if;
if pc = 56032 then
	inst <= x"03DC0070";
end if;
if pc = 56036 then
	inst <= x"037E000C";
end if;
if pc = 56040 then
	inst <= x"C57DFFFC";
end if;
if pc = 56044 then
	inst <= x"820042A4";
end if;
if pc = 56048 then
	inst <= x"07DC0070";
end if;
if pc = 56052 then
	inst <= x"8200DAF8";
end if;
if pc = 56056 then
	inst <= x"8200DAFC";
end if;
if pc = 56060 then
	inst <= x"8200DB00";
end if;
if pc = 56064 then
	inst <= x"02200370";
end if;
if pc = 56068 then
	inst <= x"005A0000";
end if;
if pc = 56072 then
	inst <= x"03BA000C";
end if;
if pc = 56076 then
	inst <= x"C83C0028";
end if;
if pc = 56080 then
	inst <= x"CC240008";
end if;
if pc = 56084 then
	inst <= x"C07C0050";
end if;
if pc = 56088 then
	inst <= x"C4640004";
end if;
if pc = 56092 then
	inst <= x"C07C0024";
end if;
if pc = 56096 then
	inst <= x"C4640000";
end if;
if pc = 56100 then
	inst <= x"C07C0020";
end if;
if pc = 56104 then
	inst <= x"22860220";
end if;
if pc = 56108 then
	inst <= x"D4428000";
end if;
if pc = 56112 then
	inst <= x"02460001";
end if;
if pc = 56116 then
	inst <= x"C09C001C";
end if;
if pc = 56120 then
	inst <= x"02A80002";
end if;
if pc = 56124 then
	inst <= x"C0DC0018";
end if;
if pc = 56128 then
	inst <= x"C84C0004";
end if;
if pc = 56132 then
	inst <= x"02E00003";
end if;
if pc = 56136 then
	inst <= x"C87C0010";
end if;
if pc = 56140 then
	inst <= x"C43C0068";
end if;
if pc = 56144 then
	inst <= x"C45C006C";
end if;
if pc = 56148 then
	inst <= x"C4BC0070";
end if;
if pc = 56152 then
	inst <= x"CC5C0078";
end if;
if pc = 56156 then
	inst <= x"C17DFFFC";
end if;
if pc = 56160 then
	inst <= x"002E0000";
end if;
if pc = 56164 then
	inst <= x"40206000";
end if;
if pc = 56168 then
	inst <= x"03DC0088";
end if;
if pc = 56172 then
	inst <= x"037E000C";
end if;
if pc = 56176 then
	inst <= x"C57DFFFC";
end if;
if pc = 56180 then
	inst <= x"8200081C";
end if;
if pc = 56184 then
	inst <= x"07DC0088";
end if;
if pc = 56188 then
	inst <= x"00420000";
end if;
if pc = 56192 then
	inst <= x"C03C0048";
end if;
if pc = 56196 then
	inst <= x"C0620000";
end if;
if pc = 56200 then
	inst <= x"C45C0080";
end if;
if pc = 56204 then
	inst <= x"C17DFFFC";
end if;
if pc = 56208 then
	inst <= x"00260000";
end if;
if pc = 56212 then
	inst <= x"03DC008C";
end if;
if pc = 56216 then
	inst <= x"037E000C";
end if;
if pc = 56220 then
	inst <= x"C57DFFFC";
end if;
if pc = 56224 then
	inst <= x"8200081C";
end if;
if pc = 56228 then
	inst <= x"07DC008C";
end if;
if pc = 56232 then
	inst <= x"005A0000";
end if;
if pc = 56236 then
	inst <= x"03BA0008";
end if;
if pc = 56240 then
	inst <= x"C4240004";
end if;
if pc = 56244 then
	inst <= x"C07C0080";
end if;
if pc = 56248 then
	inst <= x"C4640000";
end if;
if pc = 56252 then
	inst <= x"C83C0008";
end if;
if pc = 56256 then
	inst <= x"CC260000";
end if;
if pc = 56260 then
	inst <= x"C85C0078";
end if;
if pc = 56264 then
	inst <= x"CC460004";
end if;
if pc = 56268 then
	inst <= x"C85C0030";
end if;
if pc = 56272 then
	inst <= x"CC460008";
end if;
if pc = 56276 then
	inst <= x"C09C0048";
end if;
if pc = 56280 then
	inst <= x"C0A80000";
end if;
if pc = 56284 then
	inst <= x"06AA0001";
end if;
if pc = 56288 then
	inst <= x"C45C0084";
end if;
if pc = 56292 then
	inst <= x"86A0DE80";
end if;
if pc = 56296 then
	inst <= x"02C000C8";
end if;
if pc = 56300 then
	inst <= x"22EA0220";
end if;
if pc = 56304 then
	inst <= x"D0ECE000";
end if;
if pc = 56308 then
	inst <= x"C10E0004";
end if;
if pc = 56312 then
	inst <= x"03200001";
end if;
if pc = 56316 then
	inst <= x"C4DC0088";
end if;
if pc = 56320 then
	inst <= x"8312DC84";
end if;
if pc = 56324 then
	inst <= x"03200002";
end if;
if pc = 56328 then
	inst <= x"8312DC48";
end if;
if pc = 56332 then
	inst <= x"C43C008C";
end if;
if pc = 56336 then
	inst <= x"C4BC0090";
end if;
if pc = 56340 then
	inst <= x"C17DFFFC";
end if;
if pc = 56344 then
	inst <= x"004E0000";
end if;
if pc = 56348 then
	inst <= x"00260000";
end if;
if pc = 56352 then
	inst <= x"03DC009C";
end if;
if pc = 56356 then
	inst <= x"037E000C";
end if;
if pc = 56360 then
	inst <= x"C57DFFFC";
end if;
if pc = 56364 then
	inst <= x"8200400C";
end if;
if pc = 56368 then
	inst <= x"07DC009C";
end if;
if pc = 56372 then
	inst <= x"C05C0090";
end if;
if pc = 56376 then
	inst <= x"22640220";
end if;
if pc = 56380 then
	inst <= x"C09C008C";
end if;
if pc = 56384 then
	inst <= x"D4286000";
end if;
if pc = 56388 then
	inst <= x"8200DC80";
end if;
if pc = 56392 then
	inst <= x"C43C008C";
end if;
if pc = 56396 then
	inst <= x"C4BC0090";
end if;
if pc = 56400 then
	inst <= x"C17DFFFC";
end if;
if pc = 56404 then
	inst <= x"004E0000";
end if;
if pc = 56408 then
	inst <= x"00260000";
end if;
if pc = 56412 then
	inst <= x"03DC009C";
end if;
if pc = 56416 then
	inst <= x"037E000C";
end if;
if pc = 56420 then
	inst <= x"C57DFFFC";
end if;
if pc = 56424 then
	inst <= x"82003E98";
end if;
if pc = 56428 then
	inst <= x"07DC009C";
end if;
if pc = 56432 then
	inst <= x"C05C0090";
end if;
if pc = 56436 then
	inst <= x"22640220";
end if;
if pc = 56440 then
	inst <= x"C09C008C";
end if;
if pc = 56444 then
	inst <= x"D4286000";
end if;
if pc = 56448 then
	inst <= x"8200DCBC";
end if;
if pc = 56452 then
	inst <= x"C43C008C";
end if;
if pc = 56456 then
	inst <= x"C4BC0090";
end if;
if pc = 56460 then
	inst <= x"C17DFFFC";
end if;
if pc = 56464 then
	inst <= x"004E0000";
end if;
if pc = 56468 then
	inst <= x"00260000";
end if;
if pc = 56472 then
	inst <= x"03DC009C";
end if;
if pc = 56476 then
	inst <= x"037E000C";
end if;
if pc = 56480 then
	inst <= x"C57DFFFC";
end if;
if pc = 56484 then
	inst <= x"82003CC4";
end if;
if pc = 56488 then
	inst <= x"07DC009C";
end if;
if pc = 56492 then
	inst <= x"C05C0090";
end if;
if pc = 56496 then
	inst <= x"22640220";
end if;
if pc = 56500 then
	inst <= x"C09C008C";
end if;
if pc = 56504 then
	inst <= x"D4286000";
end if;
if pc = 56508 then
	inst <= x"06240001";
end if;
if pc = 56512 then
	inst <= x"8620DE7C";
end if;
if pc = 56516 then
	inst <= x"22420220";
end if;
if pc = 56520 then
	inst <= x"C07C0088";
end if;
if pc = 56524 then
	inst <= x"D0464000";
end if;
if pc = 56528 then
	inst <= x"C0A40004";
end if;
if pc = 56532 then
	inst <= x"02C00001";
end if;
if pc = 56536 then
	inst <= x"82ACDD54";
end if;
if pc = 56540 then
	inst <= x"02C00002";
end if;
if pc = 56544 then
	inst <= x"82ACDD1C";
end if;
if pc = 56548 then
	inst <= x"C0BC0080";
end if;
if pc = 56552 then
	inst <= x"C43C0094";
end if;
if pc = 56556 then
	inst <= x"C17DFFFC";
end if;
if pc = 56560 then
	inst <= x"002A0000";
end if;
if pc = 56564 then
	inst <= x"03DC00A0";
end if;
if pc = 56568 then
	inst <= x"037E000C";
end if;
if pc = 56572 then
	inst <= x"C57DFFFC";
end if;
if pc = 56576 then
	inst <= x"8200400C";
end if;
if pc = 56580 then
	inst <= x"07DC00A0";
end if;
if pc = 56584 then
	inst <= x"C05C0094";
end if;
if pc = 56588 then
	inst <= x"22640220";
end if;
if pc = 56592 then
	inst <= x"C09C008C";
end if;
if pc = 56596 then
	inst <= x"D4286000";
end if;
if pc = 56600 then
	inst <= x"8200DD50";
end if;
if pc = 56604 then
	inst <= x"C0BC0080";
end if;
if pc = 56608 then
	inst <= x"C43C0094";
end if;
if pc = 56612 then
	inst <= x"C17DFFFC";
end if;
if pc = 56616 then
	inst <= x"002A0000";
end if;
if pc = 56620 then
	inst <= x"03DC00A0";
end if;
if pc = 56624 then
	inst <= x"037E000C";
end if;
if pc = 56628 then
	inst <= x"C57DFFFC";
end if;
if pc = 56632 then
	inst <= x"82003E98";
end if;
if pc = 56636 then
	inst <= x"07DC00A0";
end if;
if pc = 56640 then
	inst <= x"C05C0094";
end if;
if pc = 56644 then
	inst <= x"22640220";
end if;
if pc = 56648 then
	inst <= x"C09C008C";
end if;
if pc = 56652 then
	inst <= x"D4286000";
end if;
if pc = 56656 then
	inst <= x"8200DD88";
end if;
if pc = 56660 then
	inst <= x"C0BC0080";
end if;
if pc = 56664 then
	inst <= x"C43C0094";
end if;
if pc = 56668 then
	inst <= x"C17DFFFC";
end if;
if pc = 56672 then
	inst <= x"002A0000";
end if;
if pc = 56676 then
	inst <= x"03DC00A0";
end if;
if pc = 56680 then
	inst <= x"037E000C";
end if;
if pc = 56684 then
	inst <= x"C57DFFFC";
end if;
if pc = 56688 then
	inst <= x"82003CC4";
end if;
if pc = 56692 then
	inst <= x"07DC00A0";
end if;
if pc = 56696 then
	inst <= x"C05C0094";
end if;
if pc = 56700 then
	inst <= x"22640220";
end if;
if pc = 56704 then
	inst <= x"C09C008C";
end if;
if pc = 56708 then
	inst <= x"D4286000";
end if;
if pc = 56712 then
	inst <= x"06240001";
end if;
if pc = 56716 then
	inst <= x"8620DE78";
end if;
if pc = 56720 then
	inst <= x"22420220";
end if;
if pc = 56724 then
	inst <= x"C07C0088";
end if;
if pc = 56728 then
	inst <= x"D0464000";
end if;
if pc = 56732 then
	inst <= x"C0640004";
end if;
if pc = 56736 then
	inst <= x"02A00001";
end if;
if pc = 56740 then
	inst <= x"826ADE20";
end if;
if pc = 56744 then
	inst <= x"02A00002";
end if;
if pc = 56748 then
	inst <= x"826ADDE8";
end if;
if pc = 56752 then
	inst <= x"C07C0080";
end if;
if pc = 56756 then
	inst <= x"C43C0098";
end if;
if pc = 56760 then
	inst <= x"C17DFFFC";
end if;
if pc = 56764 then
	inst <= x"00260000";
end if;
if pc = 56768 then
	inst <= x"03DC00A4";
end if;
if pc = 56772 then
	inst <= x"037E000C";
end if;
if pc = 56776 then
	inst <= x"C57DFFFC";
end if;
if pc = 56780 then
	inst <= x"8200400C";
end if;
if pc = 56784 then
	inst <= x"07DC00A4";
end if;
if pc = 56788 then
	inst <= x"C05C0098";
end if;
if pc = 56792 then
	inst <= x"22640220";
end if;
if pc = 56796 then
	inst <= x"C09C008C";
end if;
if pc = 56800 then
	inst <= x"D4286000";
end if;
if pc = 56804 then
	inst <= x"8200DE1C";
end if;
if pc = 56808 then
	inst <= x"C07C0080";
end if;
if pc = 56812 then
	inst <= x"C43C0098";
end if;
if pc = 56816 then
	inst <= x"C17DFFFC";
end if;
if pc = 56820 then
	inst <= x"00260000";
end if;
if pc = 56824 then
	inst <= x"03DC00A4";
end if;
if pc = 56828 then
	inst <= x"037E000C";
end if;
if pc = 56832 then
	inst <= x"C57DFFFC";
end if;
if pc = 56836 then
	inst <= x"82003E98";
end if;
if pc = 56840 then
	inst <= x"07DC00A4";
end if;
if pc = 56844 then
	inst <= x"C05C0098";
end if;
if pc = 56848 then
	inst <= x"22640220";
end if;
if pc = 56852 then
	inst <= x"C09C008C";
end if;
if pc = 56856 then
	inst <= x"D4286000";
end if;
if pc = 56860 then
	inst <= x"8200DE54";
end if;
if pc = 56864 then
	inst <= x"C07C0080";
end if;
if pc = 56868 then
	inst <= x"C43C0098";
end if;
if pc = 56872 then
	inst <= x"C17DFFFC";
end if;
if pc = 56876 then
	inst <= x"00260000";
end if;
if pc = 56880 then
	inst <= x"03DC00A4";
end if;
if pc = 56884 then
	inst <= x"037E000C";
end if;
if pc = 56888 then
	inst <= x"C57DFFFC";
end if;
if pc = 56892 then
	inst <= x"82003CC4";
end if;
if pc = 56896 then
	inst <= x"07DC00A4";
end if;
if pc = 56900 then
	inst <= x"C05C0098";
end if;
if pc = 56904 then
	inst <= x"22640220";
end if;
if pc = 56908 then
	inst <= x"C09C008C";
end if;
if pc = 56912 then
	inst <= x"D4286000";
end if;
if pc = 56916 then
	inst <= x"06440001";
end if;
if pc = 56920 then
	inst <= x"C03C0084";
end if;
if pc = 56924 then
	inst <= x"C17DFFFC";
end if;
if pc = 56928 then
	inst <= x"03DC00A4";
end if;
if pc = 56932 then
	inst <= x"037E000C";
end if;
if pc = 56936 then
	inst <= x"C57DFFFC";
end if;
if pc = 56940 then
	inst <= x"820042A4";
end if;
if pc = 56944 then
	inst <= x"07DC00A4";
end if;
if pc = 56948 then
	inst <= x"8200DE78";
end if;
if pc = 56952 then
	inst <= x"8200DE7C";
end if;
if pc = 56956 then
	inst <= x"8200DE80";
end if;
if pc = 56960 then
	inst <= x"003A0000";
end if;
if pc = 56964 then
	inst <= x"03BA000C";
end if;
if pc = 56968 then
	inst <= x"C83C0028";
end if;
if pc = 56972 then
	inst <= x"CC220008";
end if;
if pc = 56976 then
	inst <= x"C05C0084";
end if;
if pc = 56980 then
	inst <= x"C4420004";
end if;
if pc = 56984 then
	inst <= x"C05C0070";
end if;
if pc = 56988 then
	inst <= x"C4420000";
end if;
if pc = 56992 then
	inst <= x"C05C006C";
end if;
if pc = 56996 then
	inst <= x"22440220";
end if;
if pc = 57000 then
	inst <= x"C07C0068";
end if;
if pc = 57004 then
	inst <= x"D4264000";
end if;
if pc = 57008 then
	inst <= x"C03C0020";
end if;
if pc = 57012 then
	inst <= x"02420002";
end if;
if pc = 57016 then
	inst <= x"C09C001C";
end if;
if pc = 57020 then
	inst <= x"02880003";
end if;
if pc = 57024 then
	inst <= x"C0BC0018";
end if;
if pc = 57028 then
	inst <= x"C84A0008";
end if;
if pc = 57032 then
	inst <= x"02A00003";
end if;
if pc = 57036 then
	inst <= x"C87C0010";
end if;
if pc = 57040 then
	inst <= x"C45C009C";
end if;
if pc = 57044 then
	inst <= x"C49C00A0";
end if;
if pc = 57048 then
	inst <= x"CC5C00A8";
end if;
if pc = 57052 then
	inst <= x"C17DFFFC";
end if;
if pc = 57056 then
	inst <= x"002A0000";
end if;
if pc = 57060 then
	inst <= x"40206000";
end if;
if pc = 57064 then
	inst <= x"03DC00B8";
end if;
if pc = 57068 then
	inst <= x"037E000C";
end if;
if pc = 57072 then
	inst <= x"C57DFFFC";
end if;
if pc = 57076 then
	inst <= x"8200081C";
end if;
if pc = 57080 then
	inst <= x"07DC00B8";
end if;
if pc = 57084 then
	inst <= x"00420000";
end if;
if pc = 57088 then
	inst <= x"C03C0048";
end if;
if pc = 57092 then
	inst <= x"C0620000";
end if;
if pc = 57096 then
	inst <= x"C45C00B0";
end if;
if pc = 57100 then
	inst <= x"C17DFFFC";
end if;
if pc = 57104 then
	inst <= x"00260000";
end if;
if pc = 57108 then
	inst <= x"03DC00BC";
end if;
if pc = 57112 then
	inst <= x"037E000C";
end if;
if pc = 57116 then
	inst <= x"C57DFFFC";
end if;
if pc = 57120 then
	inst <= x"8200081C";
end if;
if pc = 57124 then
	inst <= x"07DC00BC";
end if;
if pc = 57128 then
	inst <= x"005A0000";
end if;
if pc = 57132 then
	inst <= x"03BA0008";
end if;
if pc = 57136 then
	inst <= x"C4240004";
end if;
if pc = 57140 then
	inst <= x"C07C00B0";
end if;
if pc = 57144 then
	inst <= x"C4640000";
end if;
if pc = 57148 then
	inst <= x"C83C0008";
end if;
if pc = 57152 then
	inst <= x"CC260000";
end if;
if pc = 57156 then
	inst <= x"C83C0038";
end if;
if pc = 57160 then
	inst <= x"CC260004";
end if;
if pc = 57164 then
	inst <= x"C83C00A8";
end if;
if pc = 57168 then
	inst <= x"CC260008";
end if;
if pc = 57172 then
	inst <= x"C09C0048";
end if;
if pc = 57176 then
	inst <= x"C0880000";
end if;
if pc = 57180 then
	inst <= x"06880001";
end if;
if pc = 57184 then
	inst <= x"C45C00B4";
end if;
if pc = 57188 then
	inst <= x"8680E200";
end if;
if pc = 57192 then
	inst <= x"02A000C8";
end if;
if pc = 57196 then
	inst <= x"22C80220";
end if;
if pc = 57200 then
	inst <= x"D0CAC000";
end if;
if pc = 57204 then
	inst <= x"C0EC0004";
end if;
if pc = 57208 then
	inst <= x"03000001";
end if;
if pc = 57212 then
	inst <= x"C4BC00B8";
end if;
if pc = 57216 then
	inst <= x"82F0E004";
end if;
if pc = 57220 then
	inst <= x"03000002";
end if;
if pc = 57224 then
	inst <= x"82F0DFC8";
end if;
if pc = 57228 then
	inst <= x"C43C00BC";
end if;
if pc = 57232 then
	inst <= x"C49C00C0";
end if;
if pc = 57236 then
	inst <= x"C17DFFFC";
end if;
if pc = 57240 then
	inst <= x"004C0000";
end if;
if pc = 57244 then
	inst <= x"00260000";
end if;
if pc = 57248 then
	inst <= x"03DC00CC";
end if;
if pc = 57252 then
	inst <= x"037E000C";
end if;
if pc = 57256 then
	inst <= x"C57DFFFC";
end if;
if pc = 57260 then
	inst <= x"8200400C";
end if;
if pc = 57264 then
	inst <= x"07DC00CC";
end if;
if pc = 57268 then
	inst <= x"C05C00C0";
end if;
if pc = 57272 then
	inst <= x"22640220";
end if;
if pc = 57276 then
	inst <= x"C09C00BC";
end if;
if pc = 57280 then
	inst <= x"D4286000";
end if;
if pc = 57284 then
	inst <= x"8200E000";
end if;
if pc = 57288 then
	inst <= x"C43C00BC";
end if;
if pc = 57292 then
	inst <= x"C49C00C0";
end if;
if pc = 57296 then
	inst <= x"C17DFFFC";
end if;
if pc = 57300 then
	inst <= x"004C0000";
end if;
if pc = 57304 then
	inst <= x"00260000";
end if;
if pc = 57308 then
	inst <= x"03DC00CC";
end if;
if pc = 57312 then
	inst <= x"037E000C";
end if;
if pc = 57316 then
	inst <= x"C57DFFFC";
end if;
if pc = 57320 then
	inst <= x"82003E98";
end if;
if pc = 57324 then
	inst <= x"07DC00CC";
end if;
if pc = 57328 then
	inst <= x"C05C00C0";
end if;
if pc = 57332 then
	inst <= x"22640220";
end if;
if pc = 57336 then
	inst <= x"C09C00BC";
end if;
if pc = 57340 then
	inst <= x"D4286000";
end if;
if pc = 57344 then
	inst <= x"8200E03C";
end if;
if pc = 57348 then
	inst <= x"C43C00BC";
end if;
if pc = 57352 then
	inst <= x"C49C00C0";
end if;
if pc = 57356 then
	inst <= x"C17DFFFC";
end if;
if pc = 57360 then
	inst <= x"004C0000";
end if;
if pc = 57364 then
	inst <= x"00260000";
end if;
if pc = 57368 then
	inst <= x"03DC00CC";
end if;
if pc = 57372 then
	inst <= x"037E000C";
end if;
if pc = 57376 then
	inst <= x"C57DFFFC";
end if;
if pc = 57380 then
	inst <= x"82003CC4";
end if;
if pc = 57384 then
	inst <= x"07DC00CC";
end if;
if pc = 57388 then
	inst <= x"C05C00C0";
end if;
if pc = 57392 then
	inst <= x"22640220";
end if;
if pc = 57396 then
	inst <= x"C09C00BC";
end if;
if pc = 57400 then
	inst <= x"D4286000";
end if;
if pc = 57404 then
	inst <= x"06240001";
end if;
if pc = 57408 then
	inst <= x"8620E1FC";
end if;
if pc = 57412 then
	inst <= x"22420220";
end if;
if pc = 57416 then
	inst <= x"C07C00B8";
end if;
if pc = 57420 then
	inst <= x"D0464000";
end if;
if pc = 57424 then
	inst <= x"C0A40004";
end if;
if pc = 57428 then
	inst <= x"02C00001";
end if;
if pc = 57432 then
	inst <= x"82ACE0D4";
end if;
if pc = 57436 then
	inst <= x"02C00002";
end if;
if pc = 57440 then
	inst <= x"82ACE09C";
end if;
if pc = 57444 then
	inst <= x"C0BC00B0";
end if;
if pc = 57448 then
	inst <= x"C43C00C4";
end if;
if pc = 57452 then
	inst <= x"C17DFFFC";
end if;
if pc = 57456 then
	inst <= x"002A0000";
end if;
if pc = 57460 then
	inst <= x"03DC00D0";
end if;
if pc = 57464 then
	inst <= x"037E000C";
end if;
if pc = 57468 then
	inst <= x"C57DFFFC";
end if;
if pc = 57472 then
	inst <= x"8200400C";
end if;
if pc = 57476 then
	inst <= x"07DC00D0";
end if;
if pc = 57480 then
	inst <= x"C05C00C4";
end if;
if pc = 57484 then
	inst <= x"22640220";
end if;
if pc = 57488 then
	inst <= x"C09C00BC";
end if;
if pc = 57492 then
	inst <= x"D4286000";
end if;
if pc = 57496 then
	inst <= x"8200E0D0";
end if;
if pc = 57500 then
	inst <= x"C0BC00B0";
end if;
if pc = 57504 then
	inst <= x"C43C00C4";
end if;
if pc = 57508 then
	inst <= x"C17DFFFC";
end if;
if pc = 57512 then
	inst <= x"002A0000";
end if;
if pc = 57516 then
	inst <= x"03DC00D0";
end if;
if pc = 57520 then
	inst <= x"037E000C";
end if;
if pc = 57524 then
	inst <= x"C57DFFFC";
end if;
if pc = 57528 then
	inst <= x"82003E98";
end if;
if pc = 57532 then
	inst <= x"07DC00D0";
end if;
if pc = 57536 then
	inst <= x"C05C00C4";
end if;
if pc = 57540 then
	inst <= x"22640220";
end if;
if pc = 57544 then
	inst <= x"C09C00BC";
end if;
if pc = 57548 then
	inst <= x"D4286000";
end if;
if pc = 57552 then
	inst <= x"8200E108";
end if;
if pc = 57556 then
	inst <= x"C0BC00B0";
end if;
if pc = 57560 then
	inst <= x"C43C00C4";
end if;
if pc = 57564 then
	inst <= x"C17DFFFC";
end if;
if pc = 57568 then
	inst <= x"002A0000";
end if;
if pc = 57572 then
	inst <= x"03DC00D0";
end if;
if pc = 57576 then
	inst <= x"037E000C";
end if;
if pc = 57580 then
	inst <= x"C57DFFFC";
end if;
if pc = 57584 then
	inst <= x"82003CC4";
end if;
if pc = 57588 then
	inst <= x"07DC00D0";
end if;
if pc = 57592 then
	inst <= x"C05C00C4";
end if;
if pc = 57596 then
	inst <= x"22640220";
end if;
if pc = 57600 then
	inst <= x"C09C00BC";
end if;
if pc = 57604 then
	inst <= x"D4286000";
end if;
if pc = 57608 then
	inst <= x"06240001";
end if;
if pc = 57612 then
	inst <= x"8620E1F8";
end if;
if pc = 57616 then
	inst <= x"22420220";
end if;
if pc = 57620 then
	inst <= x"C07C00B8";
end if;
if pc = 57624 then
	inst <= x"D0464000";
end if;
if pc = 57628 then
	inst <= x"C0640004";
end if;
if pc = 57632 then
	inst <= x"02A00001";
end if;
if pc = 57636 then
	inst <= x"826AE1A0";
end if;
if pc = 57640 then
	inst <= x"02A00002";
end if;
if pc = 57644 then
	inst <= x"826AE168";
end if;
if pc = 57648 then
	inst <= x"C07C00B0";
end if;
if pc = 57652 then
	inst <= x"C43C00C8";
end if;
if pc = 57656 then
	inst <= x"C17DFFFC";
end if;
if pc = 57660 then
	inst <= x"00260000";
end if;
if pc = 57664 then
	inst <= x"03DC00D4";
end if;
if pc = 57668 then
	inst <= x"037E000C";
end if;
if pc = 57672 then
	inst <= x"C57DFFFC";
end if;
if pc = 57676 then
	inst <= x"8200400C";
end if;
if pc = 57680 then
	inst <= x"07DC00D4";
end if;
if pc = 57684 then
	inst <= x"C05C00C8";
end if;
if pc = 57688 then
	inst <= x"22640220";
end if;
if pc = 57692 then
	inst <= x"C09C00BC";
end if;
if pc = 57696 then
	inst <= x"D4286000";
end if;
if pc = 57700 then
	inst <= x"8200E19C";
end if;
if pc = 57704 then
	inst <= x"C07C00B0";
end if;
if pc = 57708 then
	inst <= x"C43C00C8";
end if;
if pc = 57712 then
	inst <= x"C17DFFFC";
end if;
if pc = 57716 then
	inst <= x"00260000";
end if;
if pc = 57720 then
	inst <= x"03DC00D4";
end if;
if pc = 57724 then
	inst <= x"037E000C";
end if;
if pc = 57728 then
	inst <= x"C57DFFFC";
end if;
if pc = 57732 then
	inst <= x"82003E98";
end if;
if pc = 57736 then
	inst <= x"07DC00D4";
end if;
if pc = 57740 then
	inst <= x"C05C00C8";
end if;
if pc = 57744 then
	inst <= x"22640220";
end if;
if pc = 57748 then
	inst <= x"C09C00BC";
end if;
if pc = 57752 then
	inst <= x"D4286000";
end if;
if pc = 57756 then
	inst <= x"8200E1D4";
end if;
if pc = 57760 then
	inst <= x"C07C00B0";
end if;
if pc = 57764 then
	inst <= x"C43C00C8";
end if;
if pc = 57768 then
	inst <= x"C17DFFFC";
end if;
if pc = 57772 then
	inst <= x"00260000";
end if;
if pc = 57776 then
	inst <= x"03DC00D4";
end if;
if pc = 57780 then
	inst <= x"037E000C";
end if;
if pc = 57784 then
	inst <= x"C57DFFFC";
end if;
if pc = 57788 then
	inst <= x"82003CC4";
end if;
if pc = 57792 then
	inst <= x"07DC00D4";
end if;
if pc = 57796 then
	inst <= x"C05C00C8";
end if;
if pc = 57800 then
	inst <= x"22640220";
end if;
if pc = 57804 then
	inst <= x"C09C00BC";
end if;
if pc = 57808 then
	inst <= x"D4286000";
end if;
if pc = 57812 then
	inst <= x"06440001";
end if;
if pc = 57816 then
	inst <= x"C03C00B4";
end if;
if pc = 57820 then
	inst <= x"C17DFFFC";
end if;
if pc = 57824 then
	inst <= x"03DC00D4";
end if;
if pc = 57828 then
	inst <= x"037E000C";
end if;
if pc = 57832 then
	inst <= x"C57DFFFC";
end if;
if pc = 57836 then
	inst <= x"820042A4";
end if;
if pc = 57840 then
	inst <= x"07DC00D4";
end if;
if pc = 57844 then
	inst <= x"8200E1F8";
end if;
if pc = 57848 then
	inst <= x"8200E1FC";
end if;
if pc = 57852 then
	inst <= x"8200E200";
end if;
if pc = 57856 then
	inst <= x"003A0000";
end if;
if pc = 57860 then
	inst <= x"03BA000C";
end if;
if pc = 57864 then
	inst <= x"C83C0028";
end if;
if pc = 57868 then
	inst <= x"CC220008";
end if;
if pc = 57872 then
	inst <= x"C05C00B4";
end if;
if pc = 57876 then
	inst <= x"C4420004";
end if;
if pc = 57880 then
	inst <= x"C05C00A0";
end if;
if pc = 57884 then
	inst <= x"C4420000";
end if;
if pc = 57888 then
	inst <= x"C05C009C";
end if;
if pc = 57892 then
	inst <= x"22440220";
end if;
if pc = 57896 then
	inst <= x"C07C0068";
end if;
if pc = 57900 then
	inst <= x"D4264000";
end if;
if pc = 57904 then
	inst <= x"C03C0020";
end if;
if pc = 57908 then
	inst <= x"02220003";
end if;
if pc = 57912 then
	inst <= x"C05C0000";
end if;
if pc = 57916 then
	inst <= x"C4240000";
end if;
if pc = 57920 then
	inst <= x"C1FDFFFC";
end if;
if pc = 57924 then
	inst <= x"22220220";
end if;
if pc = 57928 then
	inst <= x"02220001";
end if;
if pc = 57932 then
	inst <= x"02600640";
end if;
if pc = 57936 then
	inst <= x"C0860000";
end if;
if pc = 57940 then
	inst <= x"C82000A8";
end if;
if pc = 57944 then
	inst <= x"C0A4001C";
end if;
if pc = 57948 then
	inst <= x"C84A0000";
end if;
if pc = 57952 then
	inst <= x"44224000";
end if;
if pc = 57956 then
	inst <= x"02A001D0";
end if;
if pc = 57960 then
	inst <= x"C0C40010";
end if;
if pc = 57964 then
	inst <= x"C84A0000";
end if;
if pc = 57968 then
	inst <= x"C86C0000";
end if;
if pc = 57972 then
	inst <= x"48446000";
end if;
if pc = 57976 then
	inst <= x"C86A0004";
end if;
if pc = 57980 then
	inst <= x"C88C0004";
end if;
if pc = 57984 then
	inst <= x"48668000";
end if;
if pc = 57988 then
	inst <= x"40446000";
end if;
if pc = 57992 then
	inst <= x"C86A0008";
end if;
if pc = 57996 then
	inst <= x"C88C0008";
end if;
if pc = 58000 then
	inst <= x"48668000";
end if;
if pc = 58004 then
	inst <= x"40446000";
end if;
if pc = 58008 then
	inst <= x"C8600080";
end if;
if pc = 58012 then
	inst <= x"C0C40010";
end if;
if pc = 58016 then
	inst <= x"C88C0000";
end if;
if pc = 58020 then
	inst <= x"48868000";
end if;
if pc = 58024 then
	inst <= x"48884000";
end if;
if pc = 58028 then
	inst <= x"C8AA0000";
end if;
if pc = 58032 then
	inst <= x"4488A000";
end if;
if pc = 58036 then
	inst <= x"C0C40010";
end if;
if pc = 58040 then
	inst <= x"C8AC0004";
end if;
if pc = 58044 then
	inst <= x"48A6A000";
end if;
if pc = 58048 then
	inst <= x"48AA4000";
end if;
if pc = 58052 then
	inst <= x"C8CA0004";
end if;
if pc = 58056 then
	inst <= x"44AAC000";
end if;
if pc = 58060 then
	inst <= x"C0440010";
end if;
if pc = 58064 then
	inst <= x"C8C40008";
end if;
if pc = 58068 then
	inst <= x"4866C000";
end if;
if pc = 58072 then
	inst <= x"48464000";
end if;
if pc = 58076 then
	inst <= x"C86A0008";
end if;
if pc = 58080 then
	inst <= x"44446000";
end if;
if pc = 58084 then
	inst <= x"02400003";
end if;
if pc = 58088 then
	inst <= x"40600000";
end if;
if pc = 58092 then
	inst <= x"C47C0000";
end if;
if pc = 58096 then
	inst <= x"C49C0004";
end if;
if pc = 58100 then
	inst <= x"C43C0008";
end if;
if pc = 58104 then
	inst <= x"CC3C0010";
end if;
if pc = 58108 then
	inst <= x"CC5C0018";
end if;
if pc = 58112 then
	inst <= x"CCBC0020";
end if;
if pc = 58116 then
	inst <= x"CC9C0028";
end if;
if pc = 58120 then
	inst <= x"C17DFFFC";
end if;
if pc = 58124 then
	inst <= x"00240000";
end if;
if pc = 58128 then
	inst <= x"40206000";
end if;
if pc = 58132 then
	inst <= x"03DC0038";
end if;
if pc = 58136 then
	inst <= x"037E000C";
end if;
if pc = 58140 then
	inst <= x"C57DFFFC";
end if;
if pc = 58144 then
	inst <= x"8200081C";
end if;
if pc = 58148 then
	inst <= x"07DC0038";
end if;
if pc = 58152 then
	inst <= x"00420000";
end if;
if pc = 58156 then
	inst <= x"022000C4";
end if;
if pc = 58160 then
	inst <= x"C0620000";
end if;
if pc = 58164 then
	inst <= x"C43C0030";
end if;
if pc = 58168 then
	inst <= x"C45C0034";
end if;
if pc = 58172 then
	inst <= x"C17DFFFC";
end if;
if pc = 58176 then
	inst <= x"00260000";
end if;
if pc = 58180 then
	inst <= x"03DC0040";
end if;
if pc = 58184 then
	inst <= x"037E000C";
end if;
if pc = 58188 then
	inst <= x"C57DFFFC";
end if;
if pc = 58192 then
	inst <= x"8200081C";
end if;
if pc = 58196 then
	inst <= x"07DC0040";
end if;
if pc = 58200 then
	inst <= x"005A0000";
end if;
if pc = 58204 then
	inst <= x"03BA0008";
end if;
if pc = 58208 then
	inst <= x"C4240004";
end if;
if pc = 58212 then
	inst <= x"C07C0034";
end if;
if pc = 58216 then
	inst <= x"C4640000";
end if;
if pc = 58220 then
	inst <= x"C83C0028";
end if;
if pc = 58224 then
	inst <= x"CC260000";
end if;
if pc = 58228 then
	inst <= x"C83C0020";
end if;
if pc = 58232 then
	inst <= x"CC260004";
end if;
if pc = 58236 then
	inst <= x"C83C0018";
end if;
if pc = 58240 then
	inst <= x"CC260008";
end if;
if pc = 58244 then
	inst <= x"C09C0030";
end if;
if pc = 58248 then
	inst <= x"C0880000";
end if;
if pc = 58252 then
	inst <= x"06880001";
end if;
if pc = 58256 then
	inst <= x"C45C0038";
end if;
if pc = 58260 then
	inst <= x"8680E630";
end if;
if pc = 58264 then
	inst <= x"02A000C8";
end if;
if pc = 58268 then
	inst <= x"22C80220";
end if;
if pc = 58272 then
	inst <= x"D0CAC000";
end if;
if pc = 58276 then
	inst <= x"C0EC0004";
end if;
if pc = 58280 then
	inst <= x"03000001";
end if;
if pc = 58284 then
	inst <= x"C4BC003C";
end if;
if pc = 58288 then
	inst <= x"82F0E434";
end if;
if pc = 58292 then
	inst <= x"03000002";
end if;
if pc = 58296 then
	inst <= x"82F0E3F8";
end if;
if pc = 58300 then
	inst <= x"C43C0040";
end if;
if pc = 58304 then
	inst <= x"C49C0044";
end if;
if pc = 58308 then
	inst <= x"C17DFFFC";
end if;
if pc = 58312 then
	inst <= x"004C0000";
end if;
if pc = 58316 then
	inst <= x"00260000";
end if;
if pc = 58320 then
	inst <= x"03DC0050";
end if;
if pc = 58324 then
	inst <= x"037E000C";
end if;
if pc = 58328 then
	inst <= x"C57DFFFC";
end if;
if pc = 58332 then
	inst <= x"8200400C";
end if;
if pc = 58336 then
	inst <= x"07DC0050";
end if;
if pc = 58340 then
	inst <= x"C05C0044";
end if;
if pc = 58344 then
	inst <= x"22640220";
end if;
if pc = 58348 then
	inst <= x"C09C0040";
end if;
if pc = 58352 then
	inst <= x"D4286000";
end if;
if pc = 58356 then
	inst <= x"8200E430";
end if;
if pc = 58360 then
	inst <= x"C43C0040";
end if;
if pc = 58364 then
	inst <= x"C49C0044";
end if;
if pc = 58368 then
	inst <= x"C17DFFFC";
end if;
if pc = 58372 then
	inst <= x"004C0000";
end if;
if pc = 58376 then
	inst <= x"00260000";
end if;
if pc = 58380 then
	inst <= x"03DC0050";
end if;
if pc = 58384 then
	inst <= x"037E000C";
end if;
if pc = 58388 then
	inst <= x"C57DFFFC";
end if;
if pc = 58392 then
	inst <= x"82003E98";
end if;
if pc = 58396 then
	inst <= x"07DC0050";
end if;
if pc = 58400 then
	inst <= x"C05C0044";
end if;
if pc = 58404 then
	inst <= x"22640220";
end if;
if pc = 58408 then
	inst <= x"C09C0040";
end if;
if pc = 58412 then
	inst <= x"D4286000";
end if;
if pc = 58416 then
	inst <= x"8200E46C";
end if;
if pc = 58420 then
	inst <= x"C43C0040";
end if;
if pc = 58424 then
	inst <= x"C49C0044";
end if;
if pc = 58428 then
	inst <= x"C17DFFFC";
end if;
if pc = 58432 then
	inst <= x"004C0000";
end if;
if pc = 58436 then
	inst <= x"00260000";
end if;
if pc = 58440 then
	inst <= x"03DC0050";
end if;
if pc = 58444 then
	inst <= x"037E000C";
end if;
if pc = 58448 then
	inst <= x"C57DFFFC";
end if;
if pc = 58452 then
	inst <= x"82003CC4";
end if;
if pc = 58456 then
	inst <= x"07DC0050";
end if;
if pc = 58460 then
	inst <= x"C05C0044";
end if;
if pc = 58464 then
	inst <= x"22640220";
end if;
if pc = 58468 then
	inst <= x"C09C0040";
end if;
if pc = 58472 then
	inst <= x"D4286000";
end if;
if pc = 58476 then
	inst <= x"06240001";
end if;
if pc = 58480 then
	inst <= x"8620E62C";
end if;
if pc = 58484 then
	inst <= x"22420220";
end if;
if pc = 58488 then
	inst <= x"C07C003C";
end if;
if pc = 58492 then
	inst <= x"D0464000";
end if;
if pc = 58496 then
	inst <= x"C0A40004";
end if;
if pc = 58500 then
	inst <= x"02C00001";
end if;
if pc = 58504 then
	inst <= x"82ACE504";
end if;
if pc = 58508 then
	inst <= x"02C00002";
end if;
if pc = 58512 then
	inst <= x"82ACE4CC";
end if;
if pc = 58516 then
	inst <= x"C0BC0034";
end if;
if pc = 58520 then
	inst <= x"C43C0048";
end if;
if pc = 58524 then
	inst <= x"C17DFFFC";
end if;
if pc = 58528 then
	inst <= x"002A0000";
end if;
if pc = 58532 then
	inst <= x"03DC0054";
end if;
if pc = 58536 then
	inst <= x"037E000C";
end if;
if pc = 58540 then
	inst <= x"C57DFFFC";
end if;
if pc = 58544 then
	inst <= x"8200400C";
end if;
if pc = 58548 then
	inst <= x"07DC0054";
end if;
if pc = 58552 then
	inst <= x"C05C0048";
end if;
if pc = 58556 then
	inst <= x"22640220";
end if;
if pc = 58560 then
	inst <= x"C09C0040";
end if;
if pc = 58564 then
	inst <= x"D4286000";
end if;
if pc = 58568 then
	inst <= x"8200E500";
end if;
if pc = 58572 then
	inst <= x"C0BC0034";
end if;
if pc = 58576 then
	inst <= x"C43C0048";
end if;
if pc = 58580 then
	inst <= x"C17DFFFC";
end if;
if pc = 58584 then
	inst <= x"002A0000";
end if;
if pc = 58588 then
	inst <= x"03DC0054";
end if;
if pc = 58592 then
	inst <= x"037E000C";
end if;
if pc = 58596 then
	inst <= x"C57DFFFC";
end if;
if pc = 58600 then
	inst <= x"82003E98";
end if;
if pc = 58604 then
	inst <= x"07DC0054";
end if;
if pc = 58608 then
	inst <= x"C05C0048";
end if;
if pc = 58612 then
	inst <= x"22640220";
end if;
if pc = 58616 then
	inst <= x"C09C0040";
end if;
if pc = 58620 then
	inst <= x"D4286000";
end if;
if pc = 58624 then
	inst <= x"8200E538";
end if;
if pc = 58628 then
	inst <= x"C0BC0034";
end if;
if pc = 58632 then
	inst <= x"C43C0048";
end if;
if pc = 58636 then
	inst <= x"C17DFFFC";
end if;
if pc = 58640 then
	inst <= x"002A0000";
end if;
if pc = 58644 then
	inst <= x"03DC0054";
end if;
if pc = 58648 then
	inst <= x"037E000C";
end if;
if pc = 58652 then
	inst <= x"C57DFFFC";
end if;
if pc = 58656 then
	inst <= x"82003CC4";
end if;
if pc = 58660 then
	inst <= x"07DC0054";
end if;
if pc = 58664 then
	inst <= x"C05C0048";
end if;
if pc = 58668 then
	inst <= x"22640220";
end if;
if pc = 58672 then
	inst <= x"C09C0040";
end if;
if pc = 58676 then
	inst <= x"D4286000";
end if;
if pc = 58680 then
	inst <= x"06240001";
end if;
if pc = 58684 then
	inst <= x"8620E628";
end if;
if pc = 58688 then
	inst <= x"22420220";
end if;
if pc = 58692 then
	inst <= x"C07C003C";
end if;
if pc = 58696 then
	inst <= x"D0464000";
end if;
if pc = 58700 then
	inst <= x"C0640004";
end if;
if pc = 58704 then
	inst <= x"02A00001";
end if;
if pc = 58708 then
	inst <= x"826AE5D0";
end if;
if pc = 58712 then
	inst <= x"02A00002";
end if;
if pc = 58716 then
	inst <= x"826AE598";
end if;
if pc = 58720 then
	inst <= x"C07C0034";
end if;
if pc = 58724 then
	inst <= x"C43C004C";
end if;
if pc = 58728 then
	inst <= x"C17DFFFC";
end if;
if pc = 58732 then
	inst <= x"00260000";
end if;
if pc = 58736 then
	inst <= x"03DC0058";
end if;
if pc = 58740 then
	inst <= x"037E000C";
end if;
if pc = 58744 then
	inst <= x"C57DFFFC";
end if;
if pc = 58748 then
	inst <= x"8200400C";
end if;
if pc = 58752 then
	inst <= x"07DC0058";
end if;
if pc = 58756 then
	inst <= x"C05C004C";
end if;
if pc = 58760 then
	inst <= x"22640220";
end if;
if pc = 58764 then
	inst <= x"C09C0040";
end if;
if pc = 58768 then
	inst <= x"D4286000";
end if;
if pc = 58772 then
	inst <= x"8200E5CC";
end if;
if pc = 58776 then
	inst <= x"C07C0034";
end if;
if pc = 58780 then
	inst <= x"C43C004C";
end if;
if pc = 58784 then
	inst <= x"C17DFFFC";
end if;
if pc = 58788 then
	inst <= x"00260000";
end if;
if pc = 58792 then
	inst <= x"03DC0058";
end if;
if pc = 58796 then
	inst <= x"037E000C";
end if;
if pc = 58800 then
	inst <= x"C57DFFFC";
end if;
if pc = 58804 then
	inst <= x"82003E98";
end if;
if pc = 58808 then
	inst <= x"07DC0058";
end if;
if pc = 58812 then
	inst <= x"C05C004C";
end if;
if pc = 58816 then
	inst <= x"22640220";
end if;
if pc = 58820 then
	inst <= x"C09C0040";
end if;
if pc = 58824 then
	inst <= x"D4286000";
end if;
if pc = 58828 then
	inst <= x"8200E604";
end if;
if pc = 58832 then
	inst <= x"C07C0034";
end if;
if pc = 58836 then
	inst <= x"C43C004C";
end if;
if pc = 58840 then
	inst <= x"C17DFFFC";
end if;
if pc = 58844 then
	inst <= x"00260000";
end if;
if pc = 58848 then
	inst <= x"03DC0058";
end if;
if pc = 58852 then
	inst <= x"037E000C";
end if;
if pc = 58856 then
	inst <= x"C57DFFFC";
end if;
if pc = 58860 then
	inst <= x"82003CC4";
end if;
if pc = 58864 then
	inst <= x"07DC0058";
end if;
if pc = 58868 then
	inst <= x"C05C004C";
end if;
if pc = 58872 then
	inst <= x"22640220";
end if;
if pc = 58876 then
	inst <= x"C09C0040";
end if;
if pc = 58880 then
	inst <= x"D4286000";
end if;
if pc = 58884 then
	inst <= x"06440001";
end if;
if pc = 58888 then
	inst <= x"C03C0038";
end if;
if pc = 58892 then
	inst <= x"C17DFFFC";
end if;
if pc = 58896 then
	inst <= x"03DC0058";
end if;
if pc = 58900 then
	inst <= x"037E000C";
end if;
if pc = 58904 then
	inst <= x"C57DFFFC";
end if;
if pc = 58908 then
	inst <= x"820042A4";
end if;
if pc = 58912 then
	inst <= x"07DC0058";
end if;
if pc = 58916 then
	inst <= x"8200E628";
end if;
if pc = 58920 then
	inst <= x"8200E62C";
end if;
if pc = 58924 then
	inst <= x"8200E630";
end if;
if pc = 58928 then
	inst <= x"02200370";
end if;
if pc = 58932 then
	inst <= x"005A0000";
end if;
if pc = 58936 then
	inst <= x"03BA000C";
end if;
if pc = 58940 then
	inst <= x"C83C0010";
end if;
if pc = 58944 then
	inst <= x"CC240008";
end if;
if pc = 58948 then
	inst <= x"C07C0038";
end if;
if pc = 58952 then
	inst <= x"C4640004";
end if;
if pc = 58956 then
	inst <= x"C07C0008";
end if;
if pc = 58960 then
	inst <= x"C4640000";
end if;
if pc = 58964 then
	inst <= x"C07C0004";
end if;
if pc = 58968 then
	inst <= x"22860220";
end if;
if pc = 58972 then
	inst <= x"D4428000";
end if;
if pc = 58976 then
	inst <= x"02260001";
end if;
if pc = 58980 then
	inst <= x"C05C0000";
end if;
if pc = 58984 then
	inst <= x"C4240000";
end if;
if pc = 58988 then
	inst <= x"C1FDFFFC";
end if;
if pc = 58992 then
	inst <= x"026002F8";
end if;
if pc = 58996 then
	inst <= x"C4260000";
end if;
if pc = 59000 then
	inst <= x"C4460004";
end if;
if pc = 59004 then
	inst <= x"02800300";
end if;
if pc = 59008 then
	inst <= x"22A201A0";
end if;
if pc = 59012 then
	inst <= x"C4A80000";
end if;
if pc = 59016 then
	inst <= x"224401A0";
end if;
if pc = 59020 then
	inst <= x"C4480004";
end if;
if pc = 59024 then
	inst <= x"02400308";
end if;
if pc = 59028 then
	inst <= x"C8200004";
end if;
if pc = 59032 then
	inst <= x"58420000";
end if;
if pc = 59036 then
	inst <= x"C47C0000";
end if;
if pc = 59040 then
	inst <= x"C45C0004";
end if;
if pc = 59044 then
	inst <= x"CC3C0008";
end if;
if pc = 59048 then
	inst <= x"C17DFFFC";
end if;
if pc = 59052 then
	inst <= x"40204000";
end if;
if pc = 59056 then
	inst <= x"03DC0018";
end if;
if pc = 59060 then
	inst <= x"037E000C";
end if;
if pc = 59064 then
	inst <= x"C57DFFFC";
end if;
if pc = 59068 then
	inst <= x"82000844";
end if;
if pc = 59072 then
	inst <= x"07DC0018";
end if;
if pc = 59076 then
	inst <= x"C85C0008";
end if;
if pc = 59080 then
	inst <= x"48242000";
end if;
if pc = 59084 then
	inst <= x"C03C0004";
end if;
if pc = 59088 then
	inst <= x"CC220000";
end if;
if pc = 59092 then
	inst <= x"C03C0000";
end if;
if pc = 59096 then
	inst <= x"C0420000";
end if;
if pc = 59100 then
	inst <= x"C45C0010";
end if;
if pc = 59104 then
	inst <= x"C17DFFFC";
end if;
if pc = 59108 then
	inst <= x"03DC001C";
end if;
if pc = 59112 then
	inst <= x"037E000C";
end if;
if pc = 59116 then
	inst <= x"C57DFFFC";
end if;
if pc = 59120 then
	inst <= x"8200A47C";
end if;
if pc = 59124 then
	inst <= x"07DC001C";
end if;
if pc = 59128 then
	inst <= x"00420000";
end if;
if pc = 59132 then
	inst <= x"C03C0010";
end if;
if pc = 59136 then
	inst <= x"C17DFFFC";
end if;
if pc = 59140 then
	inst <= x"03DC001C";
end if;
if pc = 59144 then
	inst <= x"037E000C";
end if;
if pc = 59148 then
	inst <= x"C57DFFFC";
end if;
if pc = 59152 then
	inst <= x"8200081C";
end if;
if pc = 59156 then
	inst <= x"07DC001C";
end if;
if pc = 59160 then
	inst <= x"C05C0000";
end if;
if pc = 59164 then
	inst <= x"C0640000";
end if;
if pc = 59168 then
	inst <= x"06660002";
end if;
if pc = 59172 then
	inst <= x"C17DFFFC";
end if;
if pc = 59176 then
	inst <= x"00460000";
end if;
if pc = 59180 then
	inst <= x"03DC001C";
end if;
if pc = 59184 then
	inst <= x"037E000C";
end if;
if pc = 59188 then
	inst <= x"C57DFFFC";
end if;
if pc = 59192 then
	inst <= x"8200A914";
end if;
if pc = 59196 then
	inst <= x"07DC001C";
end if;
if pc = 59200 then
	inst <= x"C05C0000";
end if;
if pc = 59204 then
	inst <= x"C0640000";
end if;
if pc = 59208 then
	inst <= x"C43C0014";
end if;
if pc = 59212 then
	inst <= x"C47C0018";
end if;
if pc = 59216 then
	inst <= x"C17DFFFC";
end if;
if pc = 59220 then
	inst <= x"03DC0024";
end if;
if pc = 59224 then
	inst <= x"037E000C";
end if;
if pc = 59228 then
	inst <= x"C57DFFFC";
end if;
if pc = 59232 then
	inst <= x"8200A47C";
end if;
if pc = 59236 then
	inst <= x"07DC0024";
end if;
if pc = 59240 then
	inst <= x"00420000";
end if;
if pc = 59244 then
	inst <= x"C03C0018";
end if;
if pc = 59248 then
	inst <= x"C17DFFFC";
end if;
if pc = 59252 then
	inst <= x"03DC0024";
end if;
if pc = 59256 then
	inst <= x"037E000C";
end if;
if pc = 59260 then
	inst <= x"C57DFFFC";
end if;
if pc = 59264 then
	inst <= x"8200081C";
end if;
if pc = 59268 then
	inst <= x"07DC0024";
end if;
if pc = 59272 then
	inst <= x"C05C0000";
end if;
if pc = 59276 then
	inst <= x"C0640000";
end if;
if pc = 59280 then
	inst <= x"06660002";
end if;
if pc = 59284 then
	inst <= x"C17DFFFC";
end if;
if pc = 59288 then
	inst <= x"00460000";
end if;
if pc = 59292 then
	inst <= x"03DC0024";
end if;
if pc = 59296 then
	inst <= x"037E000C";
end if;
if pc = 59300 then
	inst <= x"C57DFFFC";
end if;
if pc = 59304 then
	inst <= x"8200A914";
end if;
if pc = 59308 then
	inst <= x"07DC0024";
end if;
if pc = 59312 then
	inst <= x"C05C0000";
end if;
if pc = 59316 then
	inst <= x"C0640000";
end if;
if pc = 59320 then
	inst <= x"C43C001C";
end if;
if pc = 59324 then
	inst <= x"C47C0020";
end if;
if pc = 59328 then
	inst <= x"C17DFFFC";
end if;
if pc = 59332 then
	inst <= x"03DC002C";
end if;
if pc = 59336 then
	inst <= x"037E000C";
end if;
if pc = 59340 then
	inst <= x"C57DFFFC";
end if;
if pc = 59344 then
	inst <= x"8200A47C";
end if;
if pc = 59348 then
	inst <= x"07DC002C";
end if;
if pc = 59352 then
	inst <= x"00420000";
end if;
if pc = 59356 then
	inst <= x"C03C0020";
end if;
if pc = 59360 then
	inst <= x"C17DFFFC";
end if;
if pc = 59364 then
	inst <= x"03DC002C";
end if;
if pc = 59368 then
	inst <= x"037E000C";
end if;
if pc = 59372 then
	inst <= x"C57DFFFC";
end if;
if pc = 59376 then
	inst <= x"8200081C";
end if;
if pc = 59380 then
	inst <= x"07DC002C";
end if;
if pc = 59384 then
	inst <= x"C05C0000";
end if;
if pc = 59388 then
	inst <= x"C0640000";
end if;
if pc = 59392 then
	inst <= x"06660002";
end if;
if pc = 59396 then
	inst <= x"C17DFFFC";
end if;
if pc = 59400 then
	inst <= x"00460000";
end if;
if pc = 59404 then
	inst <= x"03DC002C";
end if;
if pc = 59408 then
	inst <= x"037E000C";
end if;
if pc = 59412 then
	inst <= x"C57DFFFC";
end if;
if pc = 59416 then
	inst <= x"8200A914";
end if;
if pc = 59420 then
	inst <= x"07DC002C";
end if;
if pc = 59424 then
	inst <= x"C43C0024";
end if;
if pc = 59428 then
	inst <= x"C17DFFFC";
end if;
if pc = 59432 then
	inst <= x"03DC0030";
end if;
if pc = 59436 then
	inst <= x"037E000C";
end if;
if pc = 59440 then
	inst <= x"C57DFFFC";
end if;
if pc = 59444 then
	inst <= x"820016D4";
end if;
if pc = 59448 then
	inst <= x"07DC0030";
end if;
if pc = 59452 then
	inst <= x"C17DFFFC";
end if;
if pc = 59456 then
	inst <= x"03DC0030";
end if;
if pc = 59460 then
	inst <= x"037E000C";
end if;
if pc = 59464 then
	inst <= x"C57DFFFC";
end if;
if pc = 59468 then
	inst <= x"82001AB8";
end if;
if pc = 59472 then
	inst <= x"07DC0030";
end if;
if pc = 59476 then
	inst <= x"02200000";
end if;
if pc = 59480 then
	inst <= x"C43C0028";
end if;
if pc = 59484 then
	inst <= x"C17DFFFC";
end if;
if pc = 59488 then
	inst <= x"03DC0034";
end if;
if pc = 59492 then
	inst <= x"037E000C";
end if;
if pc = 59496 then
	inst <= x"C57DFFFC";
end if;
if pc = 59500 then
	inst <= x"82002384";
end if;
if pc = 59504 then
	inst <= x"07DC0034";
end if;
if pc = 59508 then
	inst <= x"8220E898";
end if;
if pc = 59512 then
	inst <= x"02200001";
end if;
if pc = 59516 then
	inst <= x"C17DFFFC";
end if;
if pc = 59520 then
	inst <= x"03DC0034";
end if;
if pc = 59524 then
	inst <= x"037E000C";
end if;
if pc = 59528 then
	inst <= x"C57DFFFC";
end if;
if pc = 59532 then
	inst <= x"82002930";
end if;
if pc = 59536 then
	inst <= x"07DC0034";
end if;
if pc = 59540 then
	inst <= x"8200E8A4";
end if;
if pc = 59544 then
	inst <= x"022000C4";
end if;
if pc = 59548 then
	inst <= x"C05C0028";
end if;
if pc = 59552 then
	inst <= x"C4420000";
end if;
if pc = 59556 then
	inst <= x"C17DFFFC";
end if;
if pc = 59560 then
	inst <= x"03DC0034";
end if;
if pc = 59564 then
	inst <= x"037E000C";
end if;
if pc = 59568 then
	inst <= x"C57DFFFC";
end if;
if pc = 59572 then
	inst <= x"82000794";
end if;
if pc = 59576 then
	inst <= x"07DC0034";
end if;
if pc = 59580 then
	inst <= x"0240FFFF";
end if;
if pc = 59584 then
	inst <= x"8224E8F4";
end if;
if pc = 59588 then
	inst <= x"02400001";
end if;
if pc = 59592 then
	inst <= x"C43C002C";
end if;
if pc = 59596 then
	inst <= x"C17DFFFC";
end if;
if pc = 59600 then
	inst <= x"00240000";
end if;
if pc = 59604 then
	inst <= x"03DC0038";
end if;
if pc = 59608 then
	inst <= x"037E000C";
end if;
if pc = 59612 then
	inst <= x"C57DFFFC";
end if;
if pc = 59616 then
	inst <= x"82002A44";
end if;
if pc = 59620 then
	inst <= x"07DC0038";
end if;
if pc = 59624 then
	inst <= x"C05C002C";
end if;
if pc = 59628 then
	inst <= x"C4420000";
end if;
if pc = 59632 then
	inst <= x"8200E914";
end if;
if pc = 59636 then
	inst <= x"02200001";
end if;
if pc = 59640 then
	inst <= x"0240FFFF";
end if;
if pc = 59644 then
	inst <= x"C17DFFFC";
end if;
if pc = 59648 then
	inst <= x"03DC0038";
end if;
if pc = 59652 then
	inst <= x"037E000C";
end if;
if pc = 59656 then
	inst <= x"C57DFFFC";
end if;
if pc = 59660 then
	inst <= x"8200081C";
end if;
if pc = 59664 then
	inst <= x"07DC0038";
end if;
if pc = 59668 then
	inst <= x"C0420000";
end if;
if pc = 59672 then
	inst <= x"0260FFFF";
end if;
if pc = 59676 then
	inst <= x"8246E980";
end if;
if pc = 59680 then
	inst <= x"024001E0";
end if;
if pc = 59684 then
	inst <= x"C4240000";
end if;
if pc = 59688 then
	inst <= x"02200000";
end if;
if pc = 59692 then
	inst <= x"C45C0030";
end if;
if pc = 59696 then
	inst <= x"C17DFFFC";
end if;
if pc = 59700 then
	inst <= x"03DC003C";
end if;
if pc = 59704 then
	inst <= x"037E000C";
end if;
if pc = 59708 then
	inst <= x"C57DFFFC";
end if;
if pc = 59712 then
	inst <= x"82002A44";
end if;
if pc = 59716 then
	inst <= x"07DC003C";
end if;
if pc = 59720 then
	inst <= x"C0420000";
end if;
if pc = 59724 then
	inst <= x"0260FFFF";
end if;
if pc = 59728 then
	inst <= x"8246E97C";
end if;
if pc = 59732 then
	inst <= x"C05C0030";
end if;
if pc = 59736 then
	inst <= x"C4240004";
end if;
if pc = 59740 then
	inst <= x"02200002";
end if;
if pc = 59744 then
	inst <= x"C17DFFFC";
end if;
if pc = 59748 then
	inst <= x"03DC003C";
end if;
if pc = 59752 then
	inst <= x"037E000C";
end if;
if pc = 59756 then
	inst <= x"C57DFFFC";
end if;
if pc = 59760 then
	inst <= x"82002E74";
end if;
if pc = 59764 then
	inst <= x"07DC003C";
end if;
if pc = 59768 then
	inst <= x"8200E97C";
end if;
if pc = 59772 then
	inst <= x"8200E980";
end if;
if pc = 59776 then
	inst <= x"022002A8";
end if;
if pc = 59780 then
	inst <= x"02400000";
end if;
if pc = 59784 then
	inst <= x"C43C0034";
end if;
if pc = 59788 then
	inst <= x"C17DFFFC";
end if;
if pc = 59792 then
	inst <= x"00240000";
end if;
if pc = 59796 then
	inst <= x"03DC0040";
end if;
if pc = 59800 then
	inst <= x"037E000C";
end if;
if pc = 59804 then
	inst <= x"C57DFFFC";
end if;
if pc = 59808 then
	inst <= x"82002BEC";
end if;
if pc = 59812 then
	inst <= x"07DC0040";
end if;
if pc = 59816 then
	inst <= x"C05C0034";
end if;
if pc = 59820 then
	inst <= x"C4240000";
end if;
if pc = 59824 then
	inst <= x"02200050";
end if;
if pc = 59828 then
	inst <= x"C17DFFFC";
end if;
if pc = 59832 then
	inst <= x"03DC0040";
end if;
if pc = 59836 then
	inst <= x"037E000C";
end if;
if pc = 59840 then
	inst <= x"C57DFFFC";
end if;
if pc = 59844 then
	inst <= x"8200078C";
end if;
if pc = 59848 then
	inst <= x"07DC0040";
end if;
if pc = 59852 then
	inst <= x"02200036";
end if;
if pc = 59856 then
	inst <= x"C17DFFFC";
end if;
if pc = 59860 then
	inst <= x"03DC0040";
end if;
if pc = 59864 then
	inst <= x"037E000C";
end if;
if pc = 59868 then
	inst <= x"C57DFFFC";
end if;
if pc = 59872 then
	inst <= x"8200078C";
end if;
if pc = 59876 then
	inst <= x"07DC0040";
end if;
if pc = 59880 then
	inst <= x"0220000A";
end if;
if pc = 59884 then
	inst <= x"C17DFFFC";
end if;
if pc = 59888 then
	inst <= x"03DC0040";
end if;
if pc = 59892 then
	inst <= x"037E000C";
end if;
if pc = 59896 then
	inst <= x"C57DFFFC";
end if;
if pc = 59900 then
	inst <= x"8200078C";
end if;
if pc = 59904 then
	inst <= x"07DC0040";
end if;
if pc = 59908 then
	inst <= x"02200031";
end if;
if pc = 59912 then
	inst <= x"C17DFFFC";
end if;
if pc = 59916 then
	inst <= x"03DC0040";
end if;
if pc = 59920 then
	inst <= x"037E000C";
end if;
if pc = 59924 then
	inst <= x"C57DFFFC";
end if;
if pc = 59928 then
	inst <= x"8200078C";
end if;
if pc = 59932 then
	inst <= x"07DC0040";
end if;
if pc = 59936 then
	inst <= x"02200032";
end if;
if pc = 59940 then
	inst <= x"C17DFFFC";
end if;
if pc = 59944 then
	inst <= x"03DC0040";
end if;
if pc = 59948 then
	inst <= x"037E000C";
end if;
if pc = 59952 then
	inst <= x"C57DFFFC";
end if;
if pc = 59956 then
	inst <= x"8200078C";
end if;
if pc = 59960 then
	inst <= x"07DC0040";
end if;
if pc = 59964 then
	inst <= x"02200038";
end if;
if pc = 59968 then
	inst <= x"C17DFFFC";
end if;
if pc = 59972 then
	inst <= x"03DC0040";
end if;
if pc = 59976 then
	inst <= x"037E000C";
end if;
if pc = 59980 then
	inst <= x"C57DFFFC";
end if;
if pc = 59984 then
	inst <= x"8200078C";
end if;
if pc = 59988 then
	inst <= x"07DC0040";
end if;
if pc = 59992 then
	inst <= x"02200020";
end if;
if pc = 59996 then
	inst <= x"C17DFFFC";
end if;
if pc = 60000 then
	inst <= x"03DC0040";
end if;
if pc = 60004 then
	inst <= x"037E000C";
end if;
if pc = 60008 then
	inst <= x"C57DFFFC";
end if;
if pc = 60012 then
	inst <= x"8200078C";
end if;
if pc = 60016 then
	inst <= x"07DC0040";
end if;
if pc = 60020 then
	inst <= x"02200031";
end if;
if pc = 60024 then
	inst <= x"C17DFFFC";
end if;
if pc = 60028 then
	inst <= x"03DC0040";
end if;
if pc = 60032 then
	inst <= x"037E000C";
end if;
if pc = 60036 then
	inst <= x"C57DFFFC";
end if;
if pc = 60040 then
	inst <= x"8200078C";
end if;
if pc = 60044 then
	inst <= x"07DC0040";
end if;
if pc = 60048 then
	inst <= x"02200032";
end if;
if pc = 60052 then
	inst <= x"C17DFFFC";
end if;
if pc = 60056 then
	inst <= x"03DC0040";
end if;
if pc = 60060 then
	inst <= x"037E000C";
end if;
if pc = 60064 then
	inst <= x"C57DFFFC";
end if;
if pc = 60068 then
	inst <= x"8200078C";
end if;
if pc = 60072 then
	inst <= x"07DC0040";
end if;
if pc = 60076 then
	inst <= x"02200038";
end if;
if pc = 60080 then
	inst <= x"C17DFFFC";
end if;
if pc = 60084 then
	inst <= x"03DC0040";
end if;
if pc = 60088 then
	inst <= x"037E000C";
end if;
if pc = 60092 then
	inst <= x"C57DFFFC";
end if;
if pc = 60096 then
	inst <= x"8200078C";
end if;
if pc = 60100 then
	inst <= x"07DC0040";
end if;
if pc = 60104 then
	inst <= x"0220000A";
end if;
if pc = 60108 then
	inst <= x"C17DFFFC";
end if;
if pc = 60112 then
	inst <= x"03DC0040";
end if;
if pc = 60116 then
	inst <= x"037E000C";
end if;
if pc = 60120 then
	inst <= x"C57DFFFC";
end if;
if pc = 60124 then
	inst <= x"8200078C";
end if;
if pc = 60128 then
	inst <= x"07DC0040";
end if;
if pc = 60132 then
	inst <= x"02200032";
end if;
if pc = 60136 then
	inst <= x"C17DFFFC";
end if;
if pc = 60140 then
	inst <= x"03DC0040";
end if;
if pc = 60144 then
	inst <= x"037E000C";
end if;
if pc = 60148 then
	inst <= x"C57DFFFC";
end if;
if pc = 60152 then
	inst <= x"8200078C";
end if;
if pc = 60156 then
	inst <= x"07DC0040";
end if;
if pc = 60160 then
	inst <= x"02200035";
end if;
if pc = 60164 then
	inst <= x"C17DFFFC";
end if;
if pc = 60168 then
	inst <= x"03DC0040";
end if;
if pc = 60172 then
	inst <= x"037E000C";
end if;
if pc = 60176 then
	inst <= x"C57DFFFC";
end if;
if pc = 60180 then
	inst <= x"8200078C";
end if;
if pc = 60184 then
	inst <= x"07DC0040";
end if;
if pc = 60188 then
	inst <= x"02200035";
end if;
if pc = 60192 then
	inst <= x"C17DFFFC";
end if;
if pc = 60196 then
	inst <= x"03DC0040";
end if;
if pc = 60200 then
	inst <= x"037E000C";
end if;
if pc = 60204 then
	inst <= x"C57DFFFC";
end if;
if pc = 60208 then
	inst <= x"8200078C";
end if;
if pc = 60212 then
	inst <= x"07DC0040";
end if;
if pc = 60216 then
	inst <= x"0220000A";
end if;
if pc = 60220 then
	inst <= x"C17DFFFC";
end if;
if pc = 60224 then
	inst <= x"03DC0040";
end if;
if pc = 60228 then
	inst <= x"037E000C";
end if;
if pc = 60232 then
	inst <= x"C57DFFFC";
end if;
if pc = 60236 then
	inst <= x"8200078C";
end if;
if pc = 60240 then
	inst <= x"07DC0040";
end if;
if pc = 60244 then
	inst <= x"02200004";
end if;
if pc = 60248 then
	inst <= x"C17DFFFC";
end if;
if pc = 60252 then
	inst <= x"03DC0040";
end if;
if pc = 60256 then
	inst <= x"037E000C";
end if;
if pc = 60260 then
	inst <= x"C57DFFFC";
end if;
if pc = 60264 then
	inst <= x"8200B92C";
end if;
if pc = 60268 then
	inst <= x"07DC0040";
end if;
if pc = 60272 then
	inst <= x"02200009";
end if;
if pc = 60276 then
	inst <= x"02400000";
end if;
if pc = 60280 then
	inst <= x"02600000";
end if;
if pc = 60284 then
	inst <= x"C17DFFFC";
end if;
if pc = 60288 then
	inst <= x"03DC0040";
end if;
if pc = 60292 then
	inst <= x"037E000C";
end if;
if pc = 60296 then
	inst <= x"C57DFFFC";
end if;
if pc = 60300 then
	inst <= x"8200B574";
end if;
if pc = 60304 then
	inst <= x"07DC0040";
end if;
if pc = 60308 then
	inst <= x"02200354";
end if;
if pc = 60312 then
	inst <= x"C0420010";
end if;
if pc = 60316 then
	inst <= x"C06401DC";
end if;
if pc = 60320 then
	inst <= x"028000C4";
end if;
if pc = 60324 then
	inst <= x"C0A80000";
end if;
if pc = 60328 then
	inst <= x"06AA0001";
end if;
if pc = 60332 then
	inst <= x"C49C0038";
end if;
if pc = 60336 then
	inst <= x"C43C003C";
end if;
if pc = 60340 then
	inst <= x"C45C0040";
end if;
if pc = 60344 then
	inst <= x"86A0EE78";
end if;
if pc = 60348 then
	inst <= x"02C000C8";
end if;
if pc = 60352 then
	inst <= x"22EA0220";
end if;
if pc = 60356 then
	inst <= x"D0ECE000";
end if;
if pc = 60360 then
	inst <= x"C1060004";
end if;
if pc = 60364 then
	inst <= x"C1260000";
end if;
if pc = 60368 then
	inst <= x"C14E0004";
end if;
if pc = 60372 then
	inst <= x"02800001";
end if;
if pc = 60376 then
	inst <= x"C47C0044";
end if;
if pc = 60380 then
	inst <= x"C4DC0048";
end if;
if pc = 60384 then
	inst <= x"8348EC64";
end if;
if pc = 60388 then
	inst <= x"02800002";
end if;
if pc = 60392 then
	inst <= x"8348EC28";
end if;
if pc = 60396 then
	inst <= x"C51C004C";
end if;
if pc = 60400 then
	inst <= x"C4BC0050";
end if;
if pc = 60404 then
	inst <= x"C17DFFFC";
end if;
if pc = 60408 then
	inst <= x"004E0000";
end if;
if pc = 60412 then
	inst <= x"00320000";
end if;
if pc = 60416 then
	inst <= x"03DC005C";
end if;
if pc = 60420 then
	inst <= x"037E000C";
end if;
if pc = 60424 then
	inst <= x"C57DFFFC";
end if;
if pc = 60428 then
	inst <= x"8200400C";
end if;
if pc = 60432 then
	inst <= x"07DC005C";
end if;
if pc = 60436 then
	inst <= x"C05C0050";
end if;
if pc = 60440 then
	inst <= x"22640220";
end if;
if pc = 60444 then
	inst <= x"C09C004C";
end if;
if pc = 60448 then
	inst <= x"D4286000";
end if;
if pc = 60452 then
	inst <= x"8200EC60";
end if;
if pc = 60456 then
	inst <= x"C51C004C";
end if;
if pc = 60460 then
	inst <= x"C4BC0050";
end if;
if pc = 60464 then
	inst <= x"C17DFFFC";
end if;
if pc = 60468 then
	inst <= x"004E0000";
end if;
if pc = 60472 then
	inst <= x"00320000";
end if;
if pc = 60476 then
	inst <= x"03DC005C";
end if;
if pc = 60480 then
	inst <= x"037E000C";
end if;
if pc = 60484 then
	inst <= x"C57DFFFC";
end if;
if pc = 60488 then
	inst <= x"82003E98";
end if;
if pc = 60492 then
	inst <= x"07DC005C";
end if;
if pc = 60496 then
	inst <= x"C05C0050";
end if;
if pc = 60500 then
	inst <= x"22640220";
end if;
if pc = 60504 then
	inst <= x"C09C004C";
end if;
if pc = 60508 then
	inst <= x"D4286000";
end if;
if pc = 60512 then
	inst <= x"8200EC9C";
end if;
if pc = 60516 then
	inst <= x"C51C004C";
end if;
if pc = 60520 then
	inst <= x"C4BC0050";
end if;
if pc = 60524 then
	inst <= x"C17DFFFC";
end if;
if pc = 60528 then
	inst <= x"004E0000";
end if;
if pc = 60532 then
	inst <= x"00320000";
end if;
if pc = 60536 then
	inst <= x"03DC005C";
end if;
if pc = 60540 then
	inst <= x"037E000C";
end if;
if pc = 60544 then
	inst <= x"C57DFFFC";
end if;
if pc = 60548 then
	inst <= x"82003CC4";
end if;
if pc = 60552 then
	inst <= x"07DC005C";
end if;
if pc = 60556 then
	inst <= x"C05C0050";
end if;
if pc = 60560 then
	inst <= x"22640220";
end if;
if pc = 60564 then
	inst <= x"C09C004C";
end if;
if pc = 60568 then
	inst <= x"D4286000";
end if;
if pc = 60572 then
	inst <= x"06240001";
end if;
if pc = 60576 then
	inst <= x"8620EE74";
end if;
if pc = 60580 then
	inst <= x"22420220";
end if;
if pc = 60584 then
	inst <= x"C07C0048";
end if;
if pc = 60588 then
	inst <= x"D0464000";
end if;
if pc = 60592 then
	inst <= x"C09C0044";
end if;
if pc = 60596 then
	inst <= x"C0A80004";
end if;
if pc = 60600 then
	inst <= x"C0C80000";
end if;
if pc = 60604 then
	inst <= x"C0E40004";
end if;
if pc = 60608 then
	inst <= x"03000001";
end if;
if pc = 60612 then
	inst <= x"82F0ED40";
end if;
if pc = 60616 then
	inst <= x"03000002";
end if;
if pc = 60620 then
	inst <= x"82F0ED08";
end if;
if pc = 60624 then
	inst <= x"C4BC0054";
end if;
if pc = 60628 then
	inst <= x"C43C0058";
end if;
if pc = 60632 then
	inst <= x"C17DFFFC";
end if;
if pc = 60636 then
	inst <= x"002C0000";
end if;
if pc = 60640 then
	inst <= x"03DC0064";
end if;
if pc = 60644 then
	inst <= x"037E000C";
end if;
if pc = 60648 then
	inst <= x"C57DFFFC";
end if;
if pc = 60652 then
	inst <= x"8200400C";
end if;
if pc = 60656 then
	inst <= x"07DC0064";
end if;
if pc = 60660 then
	inst <= x"C05C0058";
end if;
if pc = 60664 then
	inst <= x"22640220";
end if;
if pc = 60668 then
	inst <= x"C09C0054";
end if;
if pc = 60672 then
	inst <= x"D4286000";
end if;
if pc = 60676 then
	inst <= x"8200ED3C";
end if;
if pc = 60680 then
	inst <= x"C4BC0054";
end if;
if pc = 60684 then
	inst <= x"C43C0058";
end if;
if pc = 60688 then
	inst <= x"C17DFFFC";
end if;
if pc = 60692 then
	inst <= x"002C0000";
end if;
if pc = 60696 then
	inst <= x"03DC0064";
end if;
if pc = 60700 then
	inst <= x"037E000C";
end if;
if pc = 60704 then
	inst <= x"C57DFFFC";
end if;
if pc = 60708 then
	inst <= x"82003E98";
end if;
if pc = 60712 then
	inst <= x"07DC0064";
end if;
if pc = 60716 then
	inst <= x"C05C0058";
end if;
if pc = 60720 then
	inst <= x"22640220";
end if;
if pc = 60724 then
	inst <= x"C09C0054";
end if;
if pc = 60728 then
	inst <= x"D4286000";
end if;
if pc = 60732 then
	inst <= x"8200ED74";
end if;
if pc = 60736 then
	inst <= x"C4BC0054";
end if;
if pc = 60740 then
	inst <= x"C43C0058";
end if;
if pc = 60744 then
	inst <= x"C17DFFFC";
end if;
if pc = 60748 then
	inst <= x"002C0000";
end if;
if pc = 60752 then
	inst <= x"03DC0064";
end if;
if pc = 60756 then
	inst <= x"037E000C";
end if;
if pc = 60760 then
	inst <= x"C57DFFFC";
end if;
if pc = 60764 then
	inst <= x"82003CC4";
end if;
if pc = 60768 then
	inst <= x"07DC0064";
end if;
if pc = 60772 then
	inst <= x"C05C0058";
end if;
if pc = 60776 then
	inst <= x"22640220";
end if;
if pc = 60780 then
	inst <= x"C09C0054";
end if;
if pc = 60784 then
	inst <= x"D4286000";
end if;
if pc = 60788 then
	inst <= x"06240001";
end if;
if pc = 60792 then
	inst <= x"8620EE70";
end if;
if pc = 60796 then
	inst <= x"22420220";
end if;
if pc = 60800 then
	inst <= x"C07C0048";
end if;
if pc = 60804 then
	inst <= x"D0464000";
end if;
if pc = 60808 then
	inst <= x"C07C0044";
end if;
if pc = 60812 then
	inst <= x"C0860004";
end if;
if pc = 60816 then
	inst <= x"C0A60000";
end if;
if pc = 60820 then
	inst <= x"C0C40004";
end if;
if pc = 60824 then
	inst <= x"02E00001";
end if;
if pc = 60828 then
	inst <= x"82CEEE18";
end if;
if pc = 60832 then
	inst <= x"02E00002";
end if;
if pc = 60836 then
	inst <= x"82CEEDE0";
end if;
if pc = 60840 then
	inst <= x"C49C005C";
end if;
if pc = 60844 then
	inst <= x"C43C0060";
end if;
if pc = 60848 then
	inst <= x"C17DFFFC";
end if;
if pc = 60852 then
	inst <= x"002A0000";
end if;
if pc = 60856 then
	inst <= x"03DC006C";
end if;
if pc = 60860 then
	inst <= x"037E000C";
end if;
if pc = 60864 then
	inst <= x"C57DFFFC";
end if;
if pc = 60868 then
	inst <= x"8200400C";
end if;
if pc = 60872 then
	inst <= x"07DC006C";
end if;
if pc = 60876 then
	inst <= x"C05C0060";
end if;
if pc = 60880 then
	inst <= x"22640220";
end if;
if pc = 60884 then
	inst <= x"C09C005C";
end if;
if pc = 60888 then
	inst <= x"D4286000";
end if;
if pc = 60892 then
	inst <= x"8200EE14";
end if;
if pc = 60896 then
	inst <= x"C49C005C";
end if;
if pc = 60900 then
	inst <= x"C43C0060";
end if;
if pc = 60904 then
	inst <= x"C17DFFFC";
end if;
if pc = 60908 then
	inst <= x"002A0000";
end if;
if pc = 60912 then
	inst <= x"03DC006C";
end if;
if pc = 60916 then
	inst <= x"037E000C";
end if;
if pc = 60920 then
	inst <= x"C57DFFFC";
end if;
if pc = 60924 then
	inst <= x"82003E98";
end if;
if pc = 60928 then
	inst <= x"07DC006C";
end if;
if pc = 60932 then
	inst <= x"C05C0060";
end if;
if pc = 60936 then
	inst <= x"22640220";
end if;
if pc = 60940 then
	inst <= x"C09C005C";
end if;
if pc = 60944 then
	inst <= x"D4286000";
end if;
if pc = 60948 then
	inst <= x"8200EE4C";
end if;
if pc = 60952 then
	inst <= x"C49C005C";
end if;
if pc = 60956 then
	inst <= x"C43C0060";
end if;
if pc = 60960 then
	inst <= x"C17DFFFC";
end if;
if pc = 60964 then
	inst <= x"002A0000";
end if;
if pc = 60968 then
	inst <= x"03DC006C";
end if;
if pc = 60972 then
	inst <= x"037E000C";
end if;
if pc = 60976 then
	inst <= x"C57DFFFC";
end if;
if pc = 60980 then
	inst <= x"82003CC4";
end if;
if pc = 60984 then
	inst <= x"07DC006C";
end if;
if pc = 60988 then
	inst <= x"C05C0060";
end if;
if pc = 60992 then
	inst <= x"22640220";
end if;
if pc = 60996 then
	inst <= x"C09C005C";
end if;
if pc = 61000 then
	inst <= x"D4286000";
end if;
if pc = 61004 then
	inst <= x"06440001";
end if;
if pc = 61008 then
	inst <= x"C03C0044";
end if;
if pc = 61012 then
	inst <= x"C17DFFFC";
end if;
if pc = 61016 then
	inst <= x"03DC006C";
end if;
if pc = 61020 then
	inst <= x"037E000C";
end if;
if pc = 61024 then
	inst <= x"C57DFFFC";
end if;
if pc = 61028 then
	inst <= x"820042A4";
end if;
if pc = 61032 then
	inst <= x"07DC006C";
end if;
if pc = 61036 then
	inst <= x"8200EE70";
end if;
if pc = 61040 then
	inst <= x"8200EE74";
end if;
if pc = 61044 then
	inst <= x"8200EE78";
end if;
if pc = 61048 then
	inst <= x"02400076";
end if;
if pc = 61052 then
	inst <= x"C03C0040";
end if;
if pc = 61056 then
	inst <= x"C17DFFFC";
end if;
if pc = 61060 then
	inst <= x"03DC006C";
end if;
if pc = 61064 then
	inst <= x"037E000C";
end if;
if pc = 61068 then
	inst <= x"C57DFFFC";
end if;
if pc = 61072 then
	inst <= x"8200BD10";
end if;
if pc = 61076 then
	inst <= x"07DC006C";
end if;
if pc = 61080 then
	inst <= x"C03C003C";
end if;
if pc = 61084 then
	inst <= x"C022000C";
end if;
if pc = 61088 then
	inst <= x"02400077";
end if;
if pc = 61092 then
	inst <= x"C17DFFFC";
end if;
if pc = 61096 then
	inst <= x"03DC006C";
end if;
if pc = 61100 then
	inst <= x"037E000C";
end if;
if pc = 61104 then
	inst <= x"C57DFFFC";
end if;
if pc = 61108 then
	inst <= x"8200BD10";
end if;
if pc = 61112 then
	inst <= x"07DC006C";
end if;
if pc = 61116 then
	inst <= x"02200002";
end if;
if pc = 61120 then
	inst <= x"C17DFFFC";
end if;
if pc = 61124 then
	inst <= x"03DC006C";
end if;
if pc = 61128 then
	inst <= x"037E000C";
end if;
if pc = 61132 then
	inst <= x"C57DFFFC";
end if;
if pc = 61136 then
	inst <= x"8200C714";
end if;
if pc = 61140 then
	inst <= x"07DC006C";
end if;
if pc = 61144 then
	inst <= x"02200368";
end if;
if pc = 61148 then
	inst <= x"C0420000";
end if;
if pc = 61152 then
	inst <= x"026001D0";
end if;
if pc = 61156 then
	inst <= x"C8260000";
end if;
if pc = 61160 then
	inst <= x"CC240000";
end if;
if pc = 61164 then
	inst <= x"C8260004";
end if;
if pc = 61168 then
	inst <= x"CC240004";
end if;
if pc = 61172 then
	inst <= x"C8260008";
end if;
if pc = 61176 then
	inst <= x"CC240008";
end if;
if pc = 61180 then
	inst <= x"C05C0038";
end if;
if pc = 61184 then
	inst <= x"C0640000";
end if;
if pc = 61188 then
	inst <= x"06660001";
end if;
if pc = 61192 then
	inst <= x"8660F0EC";
end if;
if pc = 61196 then
	inst <= x"028000C8";
end if;
if pc = 61200 then
	inst <= x"22A60220";
end if;
if pc = 61204 then
	inst <= x"D0A8A000";
end if;
if pc = 61208 then
	inst <= x"C0C20004";
end if;
if pc = 61212 then
	inst <= x"C0E20000";
end if;
if pc = 61216 then
	inst <= x"C10A0004";
end if;
if pc = 61220 then
	inst <= x"03200001";
end if;
if pc = 61224 then
	inst <= x"C43C0064";
end if;
if pc = 61228 then
	inst <= x"C49C0068";
end if;
if pc = 61232 then
	inst <= x"8312EFB4";
end if;
if pc = 61236 then
	inst <= x"03200002";
end if;
if pc = 61240 then
	inst <= x"8312EF78";
end if;
if pc = 61244 then
	inst <= x"C4DC006C";
end if;
if pc = 61248 then
	inst <= x"C47C0070";
end if;
if pc = 61252 then
	inst <= x"C17DFFFC";
end if;
if pc = 61256 then
	inst <= x"004A0000";
end if;
if pc = 61260 then
	inst <= x"002E0000";
end if;
if pc = 61264 then
	inst <= x"03DC007C";
end if;
if pc = 61268 then
	inst <= x"037E000C";
end if;
if pc = 61272 then
	inst <= x"C57DFFFC";
end if;
if pc = 61276 then
	inst <= x"8200400C";
end if;
if pc = 61280 then
	inst <= x"07DC007C";
end if;
if pc = 61284 then
	inst <= x"C05C0070";
end if;
if pc = 61288 then
	inst <= x"22640220";
end if;
if pc = 61292 then
	inst <= x"C09C006C";
end if;
if pc = 61296 then
	inst <= x"D4286000";
end if;
if pc = 61300 then
	inst <= x"8200EFB0";
end if;
if pc = 61304 then
	inst <= x"C4DC006C";
end if;
if pc = 61308 then
	inst <= x"C47C0070";
end if;
if pc = 61312 then
	inst <= x"C17DFFFC";
end if;
if pc = 61316 then
	inst <= x"004A0000";
end if;
if pc = 61320 then
	inst <= x"002E0000";
end if;
if pc = 61324 then
	inst <= x"03DC007C";
end if;
if pc = 61328 then
	inst <= x"037E000C";
end if;
if pc = 61332 then
	inst <= x"C57DFFFC";
end if;
if pc = 61336 then
	inst <= x"82003E98";
end if;
if pc = 61340 then
	inst <= x"07DC007C";
end if;
if pc = 61344 then
	inst <= x"C05C0070";
end if;
if pc = 61348 then
	inst <= x"22640220";
end if;
if pc = 61352 then
	inst <= x"C09C006C";
end if;
if pc = 61356 then
	inst <= x"D4286000";
end if;
if pc = 61360 then
	inst <= x"8200EFEC";
end if;
if pc = 61364 then
	inst <= x"C4DC006C";
end if;
if pc = 61368 then
	inst <= x"C47C0070";
end if;
if pc = 61372 then
	inst <= x"C17DFFFC";
end if;
if pc = 61376 then
	inst <= x"004A0000";
end if;
if pc = 61380 then
	inst <= x"002E0000";
end if;
if pc = 61384 then
	inst <= x"03DC007C";
end if;
if pc = 61388 then
	inst <= x"037E000C";
end if;
if pc = 61392 then
	inst <= x"C57DFFFC";
end if;
if pc = 61396 then
	inst <= x"82003CC4";
end if;
if pc = 61400 then
	inst <= x"07DC007C";
end if;
if pc = 61404 then
	inst <= x"C05C0070";
end if;
if pc = 61408 then
	inst <= x"22640220";
end if;
if pc = 61412 then
	inst <= x"C09C006C";
end if;
if pc = 61416 then
	inst <= x"D4286000";
end if;
if pc = 61420 then
	inst <= x"06240001";
end if;
if pc = 61424 then
	inst <= x"8620F0E8";
end if;
if pc = 61428 then
	inst <= x"22420220";
end if;
if pc = 61432 then
	inst <= x"C07C0068";
end if;
if pc = 61436 then
	inst <= x"D0464000";
end if;
if pc = 61440 then
	inst <= x"C07C0064";
end if;
if pc = 61444 then
	inst <= x"C0860004";
end if;
if pc = 61448 then
	inst <= x"C0A60000";
end if;
if pc = 61452 then
	inst <= x"C0C40004";
end if;
if pc = 61456 then
	inst <= x"02E00001";
end if;
if pc = 61460 then
	inst <= x"82CEF090";
end if;
if pc = 61464 then
	inst <= x"02E00002";
end if;
if pc = 61468 then
	inst <= x"82CEF058";
end if;
if pc = 61472 then
	inst <= x"C49C0074";
end if;
if pc = 61476 then
	inst <= x"C43C0078";
end if;
if pc = 61480 then
	inst <= x"C17DFFFC";
end if;
if pc = 61484 then
	inst <= x"002A0000";
end if;
if pc = 61488 then
	inst <= x"03DC0084";
end if;
if pc = 61492 then
	inst <= x"037E000C";
end if;
if pc = 61496 then
	inst <= x"C57DFFFC";
end if;
if pc = 61500 then
	inst <= x"8200400C";
end if;
if pc = 61504 then
	inst <= x"07DC0084";
end if;
if pc = 61508 then
	inst <= x"C05C0078";
end if;
if pc = 61512 then
	inst <= x"22640220";
end if;
if pc = 61516 then
	inst <= x"C09C0074";
end if;
if pc = 61520 then
	inst <= x"D4286000";
end if;
if pc = 61524 then
	inst <= x"8200F08C";
end if;
if pc = 61528 then
	inst <= x"C49C0074";
end if;
if pc = 61532 then
	inst <= x"C43C0078";
end if;
if pc = 61536 then
	inst <= x"C17DFFFC";
end if;
if pc = 61540 then
	inst <= x"002A0000";
end if;
if pc = 61544 then
	inst <= x"03DC0084";
end if;
if pc = 61548 then
	inst <= x"037E000C";
end if;
if pc = 61552 then
	inst <= x"C57DFFFC";
end if;
if pc = 61556 then
	inst <= x"82003E98";
end if;
if pc = 61560 then
	inst <= x"07DC0084";
end if;
if pc = 61564 then
	inst <= x"C05C0078";
end if;
if pc = 61568 then
	inst <= x"22640220";
end if;
if pc = 61572 then
	inst <= x"C09C0074";
end if;
if pc = 61576 then
	inst <= x"D4286000";
end if;
if pc = 61580 then
	inst <= x"8200F0C4";
end if;
if pc = 61584 then
	inst <= x"C49C0074";
end if;
if pc = 61588 then
	inst <= x"C43C0078";
end if;
if pc = 61592 then
	inst <= x"C17DFFFC";
end if;
if pc = 61596 then
	inst <= x"002A0000";
end if;
if pc = 61600 then
	inst <= x"03DC0084";
end if;
if pc = 61604 then
	inst <= x"037E000C";
end if;
if pc = 61608 then
	inst <= x"C57DFFFC";
end if;
if pc = 61612 then
	inst <= x"82003CC4";
end if;
if pc = 61616 then
	inst <= x"07DC0084";
end if;
if pc = 61620 then
	inst <= x"C05C0078";
end if;
if pc = 61624 then
	inst <= x"22640220";
end if;
if pc = 61628 then
	inst <= x"C09C0074";
end if;
if pc = 61632 then
	inst <= x"D4286000";
end if;
if pc = 61636 then
	inst <= x"06440001";
end if;
if pc = 61640 then
	inst <= x"C03C0064";
end if;
if pc = 61644 then
	inst <= x"C17DFFFC";
end if;
if pc = 61648 then
	inst <= x"03DC0084";
end if;
if pc = 61652 then
	inst <= x"037E000C";
end if;
if pc = 61656 then
	inst <= x"C57DFFFC";
end if;
if pc = 61660 then
	inst <= x"820042A4";
end if;
if pc = 61664 then
	inst <= x"07DC0084";
end if;
if pc = 61668 then
	inst <= x"8200F0E8";
end if;
if pc = 61672 then
	inst <= x"8200F0EC";
end if;
if pc = 61676 then
	inst <= x"C03C0038";
end if;
if pc = 61680 then
	inst <= x"C0220000";
end if;
if pc = 61684 then
	inst <= x"06220001";
end if;
if pc = 61688 then
	inst <= x"8620F17C";
end if;
if pc = 61692 then
	inst <= x"024000C8";
end if;
if pc = 61696 then
	inst <= x"22620220";
end if;
if pc = 61700 then
	inst <= x"D0446000";
end if;
if pc = 61704 then
	inst <= x"C0640008";
end if;
if pc = 61708 then
	inst <= x"02800002";
end if;
if pc = 61712 then
	inst <= x"8268F118";
end if;
if pc = 61716 then
	inst <= x"8200F178";
end if;
if pc = 61720 then
	inst <= x"C064001C";
end if;
if pc = 61724 then
	inst <= x"C8260000";
end if;
if pc = 61728 then
	inst <= x"C84000A8";
end if;
if pc = 61732 then
	inst <= x"8E24F12C";
end if;
if pc = 61736 then
	inst <= x"8200F178";
end if;
if pc = 61740 then
	inst <= x"C0640004";
end if;
if pc = 61744 then
	inst <= x"02800001";
end if;
if pc = 61748 then
	inst <= x"8268F160";
end if;
if pc = 61752 then
	inst <= x"02800002";
end if;
if pc = 61756 then
	inst <= x"8268F144";
end if;
if pc = 61760 then
	inst <= x"8200F15C";
end if;
if pc = 61764 then
	inst <= x"C17DFFFC";
end if;
if pc = 61768 then
	inst <= x"03DC0084";
end if;
if pc = 61772 then
	inst <= x"037E000C";
end if;
if pc = 61776 then
	inst <= x"C57DFFFC";
end if;
if pc = 61780 then
	inst <= x"8200E244";
end if;
if pc = 61784 then
	inst <= x"07DC0084";
end if;
if pc = 61788 then
	inst <= x"8200F178";
end if;
if pc = 61792 then
	inst <= x"C17DFFFC";
end if;
if pc = 61796 then
	inst <= x"03DC0084";
end if;
if pc = 61800 then
	inst <= x"037E000C";
end if;
if pc = 61804 then
	inst <= x"C57DFFFC";
end if;
if pc = 61808 then
	inst <= x"8200D764";
end if;
if pc = 61812 then
	inst <= x"07DC0084";
end if;
if pc = 61816 then
	inst <= x"8200F17C";
end if;
if pc = 61820 then
	inst <= x"02400000";
end if;
if pc = 61824 then
	inst <= x"02600000";
end if;
if pc = 61828 then
	inst <= x"C03C001C";
end if;
if pc = 61832 then
	inst <= x"C17DFFFC";
end if;
if pc = 61836 then
	inst <= x"03DC0084";
end if;
if pc = 61840 then
	inst <= x"037E000C";
end if;
if pc = 61844 then
	inst <= x"C57DFFFC";
end if;
if pc = 61848 then
	inst <= x"82009C08";
end if;
if pc = 61852 then
	inst <= x"07DC0084";
end if;
if pc = 61856 then
	inst <= x"02400000";
end if;
if pc = 61860 then
	inst <= x"02600002";
end if;
if pc = 61864 then
	inst <= x"C03C0000";
end if;
if pc = 61868 then
	inst <= x"C0820004";
end if;
if pc = 61872 then
	inst <= x"8608F1B8";
end if;
if pc = 61876 then
	inst <= x"C1FDFFFC";
end if;
if pc = 61880 then
	inst <= x"C0220004";
end if;
if pc = 61884 then
	inst <= x"06220001";
end if;
if pc = 61888 then
	inst <= x"C45C007C";
end if;
if pc = 61892 then
	inst <= x"8602F1CC";
end if;
if pc = 61896 then
	inst <= x"8200F1F4";
end if;
if pc = 61900 then
	inst <= x"02200001";
end if;
if pc = 61904 then
	inst <= x"C09C0024";
end if;
if pc = 61908 then
	inst <= x"C17DFFFC";
end if;
if pc = 61912 then
	inst <= x"00420000";
end if;
if pc = 61916 then
	inst <= x"00280000";
end if;
if pc = 61920 then
	inst <= x"03DC0088";
end if;
if pc = 61924 then
	inst <= x"037E000C";
end if;
if pc = 61928 then
	inst <= x"C57DFFFC";
end if;
if pc = 61932 then
	inst <= x"82009C08";
end if;
if pc = 61936 then
	inst <= x"07DC0088";
end if;
if pc = 61940 then
	inst <= x"02200000";
end if;
if pc = 61944 then
	inst <= x"C05C007C";
end if;
if pc = 61948 then
	inst <= x"C07C0014";
end if;
if pc = 61952 then
	inst <= x"C09C001C";
end if;
if pc = 61956 then
	inst <= x"C0BC0024";
end if;
if pc = 61960 then
	inst <= x"C17DFFFC";
end if;
if pc = 61964 then
	inst <= x"03DC0088";
end if;
if pc = 61968 then
	inst <= x"037E000C";
end if;
if pc = 61972 then
	inst <= x"C57DFFFC";
end if;
if pc = 61976 then
	inst <= x"82009C7C";
end if;
if pc = 61980 then
	inst <= x"07DC0088";
end if;
if pc = 61984 then
	inst <= x"02200001";
end if;
if pc = 61988 then
	inst <= x"02A00004";
end if;
if pc = 61992 then
	inst <= x"C05C001C";
end if;
if pc = 61996 then
	inst <= x"C07C0024";
end if;
if pc = 62000 then
	inst <= x"C09C0014";
end if;
if pc = 62004 then
	inst <= x"C17DFFFC";
end if;
if pc = 62008 then
	inst <= x"03DC0088";
end if;
if pc = 62012 then
	inst <= x"037E000C";
end if;
if pc = 62016 then
	inst <= x"C57DFFFC";
end if;
if pc = 62020 then
	inst <= x"8200A164";
end if;
if pc = 62024 then
	inst <= x"07DC0088";
end if;
if pc = 62028 then
	inst <= x"C1FDFFFC";
end if;
if pc = 62032 then
	inst <= x"03DC0004";
end if;
if pc = 62036 then
	inst <= x"037E000C";
end if;
if pc = 62040 then
	inst <= x"C57DFFFC";
end if;
if pc = 62044 then
	inst <= x"82000644";
end if;
if pc = 62048 then
	inst <= x"07DC0004";
end if;
if pc = 62052 then
	inst <= x"02200080";
end if;
if pc = 62056 then
	inst <= x"02400080";
end if;
if pc = 62060 then
	inst <= x"C17DFFFC";
end if;
if pc = 62064 then
	inst <= x"03DC0008";
end if;
if pc = 62068 then
	inst <= x"037E000C";
end if;
if pc = 62072 then
	inst <= x"C57DFFFC";
end if;
if pc = 62076 then
	inst <= x"8200E670";
end if;
if pc = 62080 then
	inst <= x"07DC0008";
end if;
if pc = 62084 then
	inst <= x"02200000";
end if;
if pc = 62088 then
	inst <= x"8001E000";
end if;
if pc > 62088 then
	inst <= x"FFFFFFFF";
end if;
          -- load from SRAM
          -- send to core
--          if pc > 1 then
--            --debug write 0 s1
--            inst <= x"FFFFFFFF";
--          end if;
--          if pc = 0 then
--            --read s1
--            inst <= x"E0200000";
--          end if;
--          if pc = 1 then
--            --write s1
--            inst <= x"E2200000";
--            waitwrite <= x"20000";
--          end if;
          --inst_sram_addr <= pc(19 downto 0);
          --if inst_sram_request_finished = '1' then
          --  inst <= inst_sram_getvalue;
          --end if;
          --if (inst_fetched = '1') and (inst_sram_getvalue(31 downto 20) = x"FFD") then
          --  waitwrite <= x"20000";
          --  inst_sram_request <= '0';
          --else
          --  inst_sram_request <= '1';
          --end if;
        else
          inst <= x"FFFFFFFF";
        end if;
      end if;
    end if;
  end process;
end fetch_test;

