-- Fetch.vhd
-- Read code from SRAM (Not yet)
-- send back to core.vhd

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity fetch is
  Port (
    clk : in std_logic;
    load_signal : in std_logic := '0';
    pc : in std_logic_vector(31 downto 0);
    inst_sram_request : out std_logic;
    inst_sram_addr : out std_logic_vector(19 downto 0);
    inst_sram_getvalue : in std_logic_vector(31 downto 0);
    inst_sram_request_finished : in std_logic;
    inst_fetched : in std_logic;
    inst : out std_logic_vector(31 downto 0);
    waitwrite : in std_logic_vector(19 downto 0)
  );
end fetch;

architecture fetch_test of fetch is
begin
  fetch_main: process(clk)
  begin
    if rising_edge(clk) then
      if load_signal = '1' then
        if waitwrite = 0 then
if pc = 0 then
	inst <= x"820004E8";
end if;
if pc = 4 then
	inst <= x"00000000";
end if;
if pc = 8 then
	inst <= x"3F800000";
end if;
if pc = 12 then
	inst <= x"3FC00000";
end if;
if pc = 16 then
	inst <= x"43C80000";
end if;
if pc = 20 then
	inst <= x"40800000";
end if;
if pc = 24 then
	inst <= x"E0200000";
end if;
if pc = 28 then
	inst <= x"07DC0004";
end if;
if pc = 32 then
	inst <= x"C1FC0000";
end if;
if pc = 36 then
	inst <= x"E2200000";
end if;
if pc = 40 then
	inst <= x"07DC0004";
end if;
if pc = 44 then
	inst <= x"C1FC0000";
end if;
if pc = 48 then
	inst <= x"E0200000";
end if;
if pc = 52 then
	inst <= x"E0400000";
end if;
if pc = 56 then
	inst <= x"E0600000";
end if;
if pc = 60 then
	inst <= x"E0800000";
end if;
if pc = 64 then
	inst <= x"22221820";
end if;
if pc = 68 then
	inst <= x"22441020";
end if;
if pc = 72 then
	inst <= x"22660820";
end if;
if pc = 76 then
	inst <= x"00224000";
end if;
if pc = 80 then
	inst <= x"00226000";
end if;
if pc = 84 then
	inst <= x"00228000";
end if;
if pc = 88 then
	inst <= x"07DC0004";
end if;
if pc = 92 then
	inst <= x"C1FC0000";
end if;
if pc = 96 then
	inst <= x"E0200000";
end if;
if pc = 100 then
	inst <= x"E0400000";
end if;
if pc = 104 then
	inst <= x"E0600000";
end if;
if pc = 108 then
	inst <= x"E0800000";
end if;
if pc = 112 then
	inst <= x"22221820";
end if;
if pc = 116 then
	inst <= x"22441020";
end if;
if pc = 120 then
	inst <= x"22660820";
end if;
if pc = 124 then
	inst <= x"00224000";
end if;
if pc = 128 then
	inst <= x"00226000";
end if;
if pc = 132 then
	inst <= x"00228000";
end if;
if pc = 136 then
	inst <= x"C43C0004";
end if;
if pc = 140 then
	inst <= x"C83C0004";
end if;
if pc = 144 then
	inst <= x"07DC0004";
end if;
if pc = 148 then
	inst <= x"C1FC0000";
end if;
if pc = 152 then
	inst <= x"CC3C0004";
end if;
if pc = 156 then
	inst <= x"C03C0004";
end if;
if pc = 160 then
	inst <= x"228218A0";
end if;
if pc = 164 then
	inst <= x"226210A0";
end if;
if pc = 168 then
	inst <= x"224208A0";
end if;
if pc = 172 then
	inst <= x"E2800000";
end if;
if pc = 176 then
	inst <= x"E2600000";
end if;
if pc = 180 then
	inst <= x"E2400000";
end if;
if pc = 184 then
	inst <= x"E2200000";
end if;
if pc = 188 then
	inst <= x"07DC0004";
end if;
if pc = 192 then
	inst <= x"C1FC0000";
end if;
if pc = 196 then
	inst <= x"007A0000";
end if;
if pc = 200 then
	inst <= x"822000DC";
end if;
if pc = 204 then
	inst <= x"C45A0000";
end if;
if pc = 208 then
	inst <= x"06220001";
end if;
if pc = 212 then
	inst <= x"03BA0004";
end if;
if pc = 216 then
	inst <= x"820000C8";
end if;
if pc = 220 then
	inst <= x"00260000";
end if;
if pc = 224 then
	inst <= x"07DC0004";
end if;
if pc = 228 then
	inst <= x"C1FC0000";
end if;
if pc = 232 then
	inst <= x"5F375A86";
end if;
if pc = 236 then
	inst <= x"3F000000";
end if;
if pc = 240 then
	inst <= x"3FC00000";
end if;
if pc = 244 then
	inst <= x"C86000E8";
end if;
if pc = 248 then
	inst <= x"C88000EC";
end if;
if pc = 252 then
	inst <= x"C8A000F0";
end if;
if pc = 256 then
	inst <= x"CC3C0004";
end if;
if pc = 260 then
	inst <= x"C05C0004";
end if;
if pc = 264 then
	inst <= x"C06000E8";
end if;
if pc = 268 then
	inst <= x"224401A0";
end if;
if pc = 272 then
	inst <= x"04464000";
end if;
if pc = 276 then
	inst <= x"C45C0004";
end if;
if pc = 280 then
	inst <= x"C85C0004";
end if;
if pc = 284 then
	inst <= x"48828000";
end if;
if pc = 288 then
	inst <= x"48648000";
end if;
if pc = 292 then
	inst <= x"48646000";
end if;
if pc = 296 then
	inst <= x"446A6000";
end if;
if pc = 300 then
	inst <= x"48446000";
end if;
if pc = 304 then
	inst <= x"48648000";
end if;
if pc = 308 then
	inst <= x"48646000";
end if;
if pc = 312 then
	inst <= x"446A6000";
end if;
if pc = 316 then
	inst <= x"48446000";
end if;
if pc = 320 then
	inst <= x"48648000";
end if;
if pc = 324 then
	inst <= x"48646000";
end if;
if pc = 328 then
	inst <= x"446A6000";
end if;
if pc = 332 then
	inst <= x"48446000";
end if;
if pc = 336 then
	inst <= x"48224000";
end if;
if pc = 340 then
	inst <= x"07DC0004";
end if;
if pc = 344 then
	inst <= x"C1FC0000";
end if;
if pc = 348 then
	inst <= x"3F000000";
end if;
if pc = 352 then
	inst <= x"40000000";
end if;
if pc = 356 then
	inst <= x"BFF0F0F1";
end if;
if pc = 360 then
	inst <= x"4034B4B5";
end if;
if pc = 364 then
	inst <= x"CC3C0004";
end if;
if pc = 368 then
	inst <= x"C03C0004";
end if;
if pc = 372 then
	inst <= x"224217A0";
end if;
if pc = 376 then
	inst <= x"04404000";
end if;
if pc = 380 then
	inst <= x"024400FD";
end if;
if pc = 384 then
	inst <= x"22441720";
end if;
if pc = 388 then
	inst <= x"C45C0008";
end if;
if pc = 392 then
	inst <= x"C85C0008";
end if;
if pc = 396 then
	inst <= x"C060015C";
end if;
if pc = 400 then
	inst <= x"22220920";
end if;
if pc = 404 then
	inst <= x"222209A0";
end if;
if pc = 408 then
	inst <= x"00226000";
end if;
if pc = 412 then
	inst <= x"C43C0004";
end if;
if pc = 416 then
	inst <= x"C83C0004";
end if;
if pc = 420 then
	inst <= x"C8600164";
end if;
if pc = 424 then
	inst <= x"C8800168";
end if;
if pc = 428 then
	inst <= x"48626000";
end if;
if pc = 432 then
	inst <= x"40668000";
end if;
if pc = 436 then
	inst <= x"C8A00160";
end if;
if pc = 440 then
	inst <= x"48826000";
end if;
if pc = 444 then
	inst <= x"448A8000";
end if;
if pc = 448 then
	inst <= x"48668000";
end if;
if pc = 452 then
	inst <= x"48826000";
end if;
if pc = 456 then
	inst <= x"448A8000";
end if;
if pc = 460 then
	inst <= x"48668000";
end if;
if pc = 464 then
	inst <= x"48826000";
end if;
if pc = 468 then
	inst <= x"448A8000";
end if;
if pc = 472 then
	inst <= x"48668000";
end if;
if pc = 476 then
	inst <= x"48246000";
end if;
if pc = 480 then
	inst <= x"07DC0004";
end if;
if pc = 484 then
	inst <= x"C1FC0000";
end if;
if pc = 488 then
	inst <= x"BF800000";
end if;
if pc = 492 then
	inst <= x"CC3C0000";
end if;
if pc = 496 then
	inst <= x"C03C0000";
end if;
if pc = 500 then
	inst <= x"22420120";
end if;
if pc = 504 then
	inst <= x"224418A0";
end if;
if pc = 508 then
	inst <= x"02600096";
end if;
if pc = 512 then
	inst <= x"8664027C";
end if;
if pc = 516 then
	inst <= x"8264027C";
end if;
if pc = 520 then
	inst <= x"0260007E";
end if;
if pc = 524 then
	inst <= x"86460230";
end if;
if pc = 528 then
	inst <= x"82460230";
end if;
if pc = 532 then
	inst <= x"02800096";
end if;
if pc = 536 then
	inst <= x"04884000";
end if;
if pc = 540 then
	inst <= x"206280A0";
end if;
if pc = 544 then
	inst <= x"04404000";
end if;
if pc = 548 then
	inst <= x"02840096";
end if;
if pc = 552 then
	inst <= x"20668020";
end if;
if pc = 556 then
	inst <= x"82000234";
end if;
if pc = 560 then
	inst <= x"02600000";
end if;
if pc = 564 then
	inst <= x"C45C0004";
end if;
if pc = 568 then
	inst <= x"C47C0008";
end if;
if pc = 572 then
	inst <= x"C85C0004";
end if;
if pc = 576 then
	inst <= x"C87C0008";
end if;
if pc = 580 then
	inst <= x"44404000";
end if;
if pc = 584 then
	inst <= x"CC5C0004";
end if;
if pc = 588 then
	inst <= x"C05C0000";
end if;
if pc = 592 then
	inst <= x"86460278";
end if;
if pc = 596 then
	inst <= x"82460278";
end if;
if pc = 600 then
	inst <= x"8E600268";
end if;
if pc = 604 then
	inst <= x"40206000";
end if;
if pc = 608 then
	inst <= x"07DC0004";
end if;
if pc = 612 then
	inst <= x"C1FC0000";
end if;
if pc = 616 then
	inst <= x"C84001E8";
end if;
if pc = 620 then
	inst <= x"40264000";
end if;
if pc = 624 then
	inst <= x"07DC0004";
end if;
if pc = 628 then
	inst <= x"C1FC0000";
end if;
if pc = 632 then
	inst <= x"40206000";
end if;
if pc = 636 then
	inst <= x"07DC0004";
end if;
if pc = 640 then
	inst <= x"C1FC0000";
end if;
if pc = 644 then
	inst <= x"40222000";
end if;
if pc = 648 then
	inst <= x"07DC0004";
end if;
if pc = 652 then
	inst <= x"C1FC0000";
end if;
if pc = 656 then
	inst <= x"03600000";
end if;
if pc = 660 then
	inst <= x"82360320";
end if;
if pc = 664 then
	inst <= x"44668000";
end if;
if pc = 668 then
	inst <= x"4066A000";
end if;
if pc = 672 then
	inst <= x"CCBC0000";
end if;
if pc = 676 then
	inst <= x"C43C0008";
end if;
if pc = 680 then
	inst <= x"CC7C0010";
end if;
if pc = 684 then
	inst <= x"CCDC0018";
end if;
if pc = 688 then
	inst <= x"CC5C0020";
end if;
if pc = 692 then
	inst <= x"C17DFFFC";
end if;
if pc = 696 then
	inst <= x"C57C002C";
end if;
if pc = 700 then
	inst <= x"03DC0030";
end if;
if pc = 704 then
	inst <= x"037E0010";
end if;
if pc = 708 then
	inst <= x"C57C0000";
end if;
if pc = 712 then
	inst <= x"03DC0004";
end if;
if pc = 716 then
	inst <= x"82000284";
end if;
if pc = 720 then
	inst <= x"07DC0030";
end if;
if pc = 724 then
	inst <= x"C17C002C";
end if;
if pc = 728 then
	inst <= x"C57DFFFC";
end if;
if pc = 732 then
	inst <= x"C85C0020";
end if;
if pc = 736 then
	inst <= x"48224000";
end if;
if pc = 740 then
	inst <= x"C8DC0018";
end if;
if pc = 744 then
	inst <= x"4042C000";
end if;
if pc = 748 then
	inst <= x"C83C0010";
end if;
if pc = 752 then
	inst <= x"48622000";
end if;
if pc = 756 then
	inst <= x"48844000";
end if;
if pc = 760 then
	inst <= x"03600014";
end if;
if pc = 764 then
	inst <= x"C8B60000";
end if;
if pc = 768 then
	inst <= x"40E68000";
end if;
if pc = 772 then
	inst <= x"8EAE0318";
end if;
if pc = 776 then
	inst <= x"C03C0008";
end if;
if pc = 780 then
	inst <= x"06220001";
end if;
if pc = 784 then
	inst <= x"C8BC0000";
end if;
if pc = 788 then
	inst <= x"82000290";
end if;
if pc = 792 then
	inst <= x"02200031";
end if;
if pc = 796 then
	inst <= x"82000024";
end if;
if pc = 800 then
	inst <= x"02200030";
end if;
if pc = 804 then
	inst <= x"82000024";
end if;
if pc = 808 then
	inst <= x"02600190";
end if;
if pc = 812 then
	inst <= x"86260338";
end if;
if pc = 816 then
	inst <= x"07DC0004";
end if;
if pc = 820 then
	inst <= x"C1FC0000";
end if;
if pc = 824 then
	inst <= x"58220000";
end if;
if pc = 828 then
	inst <= x"C43C0000";
end if;
if pc = 832 then
	inst <= x"C45C0004";
end if;
if pc = 836 then
	inst <= x"C17DFFFC";
end if;
if pc = 840 then
	inst <= x"C57C000C";
end if;
if pc = 844 then
	inst <= x"03DC0010";
end if;
if pc = 848 then
	inst <= x"037E0010";
end if;
if pc = 852 then
	inst <= x"C57C0000";
end if;
if pc = 856 then
	inst <= x"03DC0004";
end if;
if pc = 860 then
	inst <= x"82000284";
end if;
if pc = 864 then
	inst <= x"07DC0010";
end if;
if pc = 868 then
	inst <= x"C17C000C";
end if;
if pc = 872 then
	inst <= x"C57DFFFC";
end if;
if pc = 876 then
	inst <= x"03600010";
end if;
if pc = 880 then
	inst <= x"C8560000";
end if;
if pc = 884 then
	inst <= x"CC5C0008";
end if;
if pc = 888 then
	inst <= x"CC3C0010";
end if;
if pc = 892 then
	inst <= x"C17DFFFC";
end if;
if pc = 896 then
	inst <= x"40204000";
end if;
if pc = 900 then
	inst <= x"C57C001C";
end if;
if pc = 904 then
	inst <= x"03DC0020";
end if;
if pc = 908 then
	inst <= x"037E0010";
end if;
if pc = 912 then
	inst <= x"C57C0000";
end if;
if pc = 916 then
	inst <= x"03DC0004";
end if;
if pc = 920 then
	inst <= x"8200016C";
end if;
if pc = 924 then
	inst <= x"07DC0020";
end if;
if pc = 928 then
	inst <= x"C17C001C";
end if;
if pc = 932 then
	inst <= x"C57DFFFC";
end if;
if pc = 936 then
	inst <= x"C85C0010";
end if;
if pc = 940 then
	inst <= x"48242000";
end if;
if pc = 944 then
	inst <= x"0360000C";
end if;
if pc = 948 then
	inst <= x"C8560000";
end if;
if pc = 952 then
	inst <= x"44224000";
end if;
if pc = 956 then
	inst <= x"C03C0004";
end if;
if pc = 960 then
	inst <= x"58420000";
end if;
if pc = 964 then
	inst <= x"CC3C0018";
end if;
if pc = 968 then
	inst <= x"C17DFFFC";
end if;
if pc = 972 then
	inst <= x"40204000";
end if;
if pc = 976 then
	inst <= x"C57C0024";
end if;
if pc = 980 then
	inst <= x"03DC0028";
end if;
if pc = 984 then
	inst <= x"037E0010";
end if;
if pc = 988 then
	inst <= x"C57C0000";
end if;
if pc = 992 then
	inst <= x"03DC0004";
end if;
if pc = 996 then
	inst <= x"82000284";
end if;
if pc = 1000 then
	inst <= x"07DC0028";
end if;
if pc = 1004 then
	inst <= x"C17C0024";
end if;
if pc = 1008 then
	inst <= x"C57DFFFC";
end if;
if pc = 1012 then
	inst <= x"C85C0008";
end if;
if pc = 1016 then
	inst <= x"CC3C0020";
end if;
if pc = 1020 then
	inst <= x"C17DFFFC";
end if;
if pc = 1024 then
	inst <= x"40204000";
end if;
if pc = 1028 then
	inst <= x"C57C002C";
end if;
if pc = 1032 then
	inst <= x"03DC0030";
end if;
if pc = 1036 then
	inst <= x"037E0010";
end if;
if pc = 1040 then
	inst <= x"C57C0000";
end if;
if pc = 1044 then
	inst <= x"03DC0004";
end if;
if pc = 1048 then
	inst <= x"8200016C";
end if;
if pc = 1052 then
	inst <= x"07DC0030";
end if;
if pc = 1056 then
	inst <= x"C17C002C";
end if;
if pc = 1060 then
	inst <= x"C57DFFFC";
end if;
if pc = 1064 then
	inst <= x"C85C0020";
end if;
if pc = 1068 then
	inst <= x"48242000";
end if;
if pc = 1072 then
	inst <= x"03600008";
end if;
if pc = 1076 then
	inst <= x"C8560000";
end if;
if pc = 1080 then
	inst <= x"44C24000";
end if;
if pc = 1084 then
	inst <= x"022003E8";
end if;
if pc = 1088 then
	inst <= x"03600004";
end if;
if pc = 1092 then
	inst <= x"C8360000";
end if;
if pc = 1096 then
	inst <= x"C8BC0018";
end if;
if pc = 1100 then
	inst <= x"C17DFFFC";
end if;
if pc = 1104 then
	inst <= x"40802000";
end if;
if pc = 1108 then
	inst <= x"40602000";
end if;
if pc = 1112 then
	inst <= x"40402000";
end if;
if pc = 1116 then
	inst <= x"C57C002C";
end if;
if pc = 1120 then
	inst <= x"03DC0030";
end if;
if pc = 1124 then
	inst <= x"037E0010";
end if;
if pc = 1128 then
	inst <= x"C57C0000";
end if;
if pc = 1132 then
	inst <= x"03DC0004";
end if;
if pc = 1136 then
	inst <= x"82000290";
end if;
if pc = 1140 then
	inst <= x"07DC0030";
end if;
if pc = 1144 then
	inst <= x"C17C002C";
end if;
if pc = 1148 then
	inst <= x"C57DFFFC";
end if;
if pc = 1152 then
	inst <= x"C03C0000";
end if;
if pc = 1156 then
	inst <= x"02220001";
end if;
if pc = 1160 then
	inst <= x"C05C0004";
end if;
if pc = 1164 then
	inst <= x"82000328";
end if;
if pc = 1168 then
	inst <= x"02400190";
end if;
if pc = 1172 then
	inst <= x"862404A0";
end if;
if pc = 1176 then
	inst <= x"07DC0004";
end if;
if pc = 1180 then
	inst <= x"C1FC0000";
end if;
if pc = 1184 then
	inst <= x"02400000";
end if;
if pc = 1188 then
	inst <= x"C43C0000";
end if;
if pc = 1192 then
	inst <= x"C17DFFFC";
end if;
if pc = 1196 then
	inst <= x"01240000";
end if;
if pc = 1200 then
	inst <= x"00420000";
end if;
if pc = 1204 then
	inst <= x"00320000";
end if;
if pc = 1208 then
	inst <= x"C57C0004";
end if;
if pc = 1212 then
	inst <= x"03DC0008";
end if;
if pc = 1216 then
	inst <= x"037E0010";
end if;
if pc = 1220 then
	inst <= x"C57C0000";
end if;
if pc = 1224 then
	inst <= x"03DC0004";
end if;
if pc = 1228 then
	inst <= x"82000328";
end if;
if pc = 1232 then
	inst <= x"07DC0008";
end if;
if pc = 1236 then
	inst <= x"C17C0004";
end if;
if pc = 1240 then
	inst <= x"C57DFFFC";
end if;
if pc = 1244 then
	inst <= x"C03C0000";
end if;
if pc = 1248 then
	inst <= x"02220001";
end if;
if pc = 1252 then
	inst <= x"82000490";
end if;
if pc = 1256 then
	inst <= x"02200000";
end if;
if pc = 1260 then
	inst <= x"C17DFFFC";
end if;
if pc = 1264 then
	inst <= x"C57C0004";
end if;
if pc = 1268 then
	inst <= x"03DC0008";
end if;
if pc = 1272 then
	inst <= x"037E0010";
end if;
if pc = 1276 then
	inst <= x"C57C0000";
end if;
if pc = 1280 then
	inst <= x"03DC0004";
end if;
if pc = 1284 then
	inst <= x"82000490";
end if;
if pc = 1288 then
	inst <= x"07DC0008";
end if;
if pc = 1292 then
	inst <= x"C17C0004";
end if;
if pc = 1296 then
	inst <= x"C57DFFFC";
end if;
if pc = 1300 then
	inst <= x"8001E000";
end if;
if pc > 1300 then
	inst <= x"FFFFFFFF";
end if;
          -- load from SRAM
          -- send to core
--          if pc > 1 then
--            --debug write 0 s1
--            inst <= x"FFFFFFFF";
--          end if;
--          if pc = 0 then
--            --read s1
--            inst <= x"E0200000";
--          end if;
--          if pc = 1 then
--            --write s1
--            inst <= x"E2200000";
--            waitwrite <= x"20000";
--          end if;
          --inst_sram_addr <= pc(19 downto 0);
          --if inst_sram_request_finished = '1' then
          --  inst <= inst_sram_getvalue;
          --end if;
          --if (inst_fetched = '1') and (inst_sram_getvalue(31 downto 20) = x"FFD") then
          --  waitwrite <= x"20000";
          --  inst_sram_request <= '0';
          --else
          --  inst_sram_request <= '1';
          --end if;
        else
          inst <= x"FFFFFFFF";
        end if;
      end if;
    end if;
  end process;
end fetch_test;

